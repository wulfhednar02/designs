magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect 205776 200205 223200 203405
<< l67d44 >>
rect 222695 203080 222865 203250
rect 222235 203080 222405 203250
rect 222695 200360 222865 200530
rect 206208 201536 206378 201706
rect 222235 200360 222405 200530
rect 205813 201537 205983 201707
rect 222703 201720 222873 201890
rect 222703 201287 222873 201457
rect 222703 202153 222873 202323
rect 222703 202585 222873 202755
rect 222703 200855 222873 201025
<< l67d20 >>
rect 207285 201520 207510 201720
rect 211915 201520 212975 201720
rect 205776 201430 206095 201800
<< l68d20 >>
rect 205776 201430 206435 201800
rect 222650 200825 222925 202785
<< l68d16 >>
rect 205776 201430 206435 201800
rect 222650 200835 222925 202781
<< l68d44 >>
rect 206145 203090 206295 203240
rect 206605 203090 206755 203240
rect 207525 203090 207675 203240
rect 207985 203090 208135 203240
rect 208445 203090 208595 203240
rect 208905 203090 209055 203240
rect 209365 203090 209515 203240
rect 207065 203090 207215 203240
rect 209825 203090 209975 203240
rect 210285 203090 210435 203240
rect 211205 203090 211355 203240
rect 211665 203090 211815 203240
rect 212125 203090 212275 203240
rect 212585 203090 212735 203240
rect 213045 203090 213195 203240
rect 210745 203090 210895 203240
rect 213505 203090 213655 203240
rect 213965 203090 214115 203240
rect 214885 203090 215035 203240
rect 215345 203090 215495 203240
rect 215805 203090 215955 203240
rect 216265 203090 216415 203240
rect 216725 203090 216875 203240
rect 214425 203090 214575 203240
rect 217185 203090 217335 203240
rect 217645 203090 217795 203240
rect 218565 203090 218715 203240
rect 219025 203090 219175 203240
rect 219485 203090 219635 203240
rect 219945 203090 220095 203240
rect 220405 203090 220555 203240
rect 218105 203090 218255 203240
rect 220865 203090 221015 203240
rect 221325 203090 221475 203240
rect 221785 203090 221935 203240
rect 222245 203090 222395 203240
rect 222705 203090 222855 203240
rect 206145 200370 206295 200520
rect 206605 200370 206755 200520
rect 207525 200370 207675 200520
rect 207985 200370 208135 200520
rect 208445 200370 208595 200520
rect 208905 200370 209055 200520
rect 209365 200370 209515 200520
rect 207065 200370 207215 200520
rect 209825 200370 209975 200520
rect 210285 200370 210435 200520
rect 211205 200370 211355 200520
rect 211665 200370 211815 200520
rect 212125 200370 212275 200520
rect 212585 200370 212735 200520
rect 213045 200370 213195 200520
rect 210745 200370 210895 200520
rect 213505 200370 213655 200520
rect 213965 200370 214115 200520
rect 214885 200370 215035 200520
rect 215345 200370 215495 200520
rect 215805 200370 215955 200520
rect 216265 200370 216415 200520
rect 216725 200370 216875 200520
rect 214425 200370 214575 200520
rect 217185 200370 217335 200520
rect 217645 200370 217795 200520
rect 218565 200370 218715 200520
rect 219025 200370 219175 200520
rect 219485 200370 219635 200520
rect 219945 200370 220095 200520
rect 220405 200370 220555 200520
rect 218105 200370 218255 200520
rect 220865 200370 221015 200520
rect 221325 200370 221475 200520
rect 221785 200370 221935 200520
rect 222245 200370 222395 200520
rect 222705 200370 222855 200520
<< l69d20 >>
rect 205990 202925 223010 203405
rect 205990 200205 223010 200685
<< l69d16 >>
rect 205990 202925 223010 203405
rect 205990 200205 223010 200685
<< labels >>
rlabel l68d5 206098 201634 206098 201634 0 IN
rlabel l68d5 222797 202697 222797 202697 0 OUT
rlabel l68d5 222787 200917 222787 200917 0 OUT
rlabel l68d5 222791 201805 222791 201805 0 OUT
rlabel l69d5 206178 200438 206178 200438 0 VSS
rlabel l69d5 222820 200459 222820 200459 0 VSS
rlabel l69d5 214450 200470 214450 200470 0 VSS
rlabel l69d5 209714 200459 209714 200459 0 VSS
rlabel l69d5 219055 200492 219055 200492 0 VSS
rlabel l69d5 206298 203177 206298 203177 0 VDD
rlabel l69d5 222755 203199 222755 203199 0 VDD
rlabel l69d5 214439 203188 214439 203188 0 VDD
rlabel l69d5 209757 203177 209757 203177 0 VDD
rlabel l69d5 219153 203188 219153 203188 0 VDD
use sky130_fd_sc_hd__buf_16 sky130_fd_sc_hd__buf_16_1
timestamp 1698899266
transform 1 0 212890 0 1 200445
box -190 -240 10310 2960
use sky130_fd_sc_hd__buf_8 sky130_fd_sc_hd__buf_8_1
timestamp 1698899266
transform 1 0 207370 0 1 200445
box -190 -240 5710 2960
use sky130_fd_sc_hd__buf_1 sky130_fd_sc_hd__buf_1_1
timestamp 1698899266
transform 1 0 205990 0 1 200445
box -190 -240 1570 2960
<< end >>
