magic
tech sky130A
magscale 1 2
timestamp 1699066547
<< error_p >>
rect 92 518 162 546
<< xpolycontact >>
rect 92 518 162 954
rect 92 40 162 476
<< ppolyres >>
rect 92 476 162 518
<< viali >>
rect 110 901 144 935
rect 110 829 144 863
rect 110 757 144 791
rect 110 685 144 719
rect 110 613 144 647
rect 110 541 144 575
rect 110 420 144 454
rect 110 348 144 382
rect 110 276 144 310
rect 110 204 144 238
rect 110 132 144 166
rect 110 60 144 94
<< metal1 >>
rect 102 935 152 948
rect 102 901 110 935
rect 144 901 152 935
rect 102 863 152 901
rect 102 829 110 863
rect 144 829 152 863
rect 102 791 152 829
rect 102 757 110 791
rect 144 757 152 791
rect 102 719 152 757
rect 102 685 110 719
rect 144 685 152 719
rect 102 647 152 685
rect 102 613 110 647
rect 144 613 152 647
rect 102 575 152 613
rect 102 541 110 575
rect 144 541 152 575
rect 102 527 152 541
rect 102 454 152 467
rect 102 420 110 454
rect 144 420 152 454
rect 102 382 152 420
rect 102 348 110 382
rect 144 348 152 382
rect 102 310 152 348
rect 102 276 110 310
rect 144 276 152 310
rect 102 238 152 276
rect 102 204 110 238
rect 144 204 152 238
rect 102 166 152 204
rect 102 132 110 166
rect 144 132 152 166
rect 102 94 152 132
rect 102 60 110 94
rect 144 60 152 94
rect 102 46 152 60
<< end >>
