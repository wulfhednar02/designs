magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< nwell >>
rect 0 309 1180 630
<< pwell >>
rect 39 69 1065 251
rect 68 31 102 69
<< scnmos >>
rect 117 95 147 225
rect 201 95 231 225
rect 285 95 315 225
rect 369 95 399 225
rect 453 95 483 225
rect 537 95 567 225
rect 621 95 651 225
rect 705 95 735 225
rect 789 95 819 225
rect 873 95 903 225
rect 957 95 987 225
<< scpmoshvt >>
rect 117 345 147 545
rect 201 345 231 545
rect 285 345 315 545
rect 369 345 399 545
rect 453 345 483 545
rect 537 345 567 545
rect 621 345 651 545
rect 705 345 735 545
rect 789 345 819 545
rect 873 345 903 545
rect 957 345 987 545
<< ndiff >>
rect 65 177 117 225
rect 65 143 73 177
rect 107 143 117 177
rect 65 95 117 143
rect 147 145 201 225
rect 147 111 157 145
rect 191 111 201 145
rect 147 95 201 111
rect 231 177 285 225
rect 231 143 241 177
rect 275 143 285 177
rect 231 95 285 143
rect 315 145 369 225
rect 315 111 325 145
rect 359 111 369 145
rect 315 95 369 111
rect 399 177 453 225
rect 399 143 409 177
rect 443 143 453 177
rect 399 95 453 143
rect 483 145 537 225
rect 483 111 493 145
rect 527 111 537 145
rect 483 95 537 111
rect 567 177 621 225
rect 567 143 577 177
rect 611 143 621 177
rect 567 95 621 143
rect 651 145 705 225
rect 651 111 661 145
rect 695 111 705 145
rect 651 95 705 111
rect 735 177 789 225
rect 735 143 745 177
rect 779 143 789 177
rect 735 95 789 143
rect 819 145 873 225
rect 819 111 829 145
rect 863 111 873 145
rect 819 95 873 111
rect 903 177 957 225
rect 903 143 913 177
rect 947 143 957 177
rect 903 95 957 143
rect 987 209 1039 225
rect 987 175 997 209
rect 1031 175 1039 209
rect 987 141 1039 175
rect 987 107 997 141
rect 1031 107 1039 141
rect 987 95 1039 107
<< pdiff >>
rect 65 527 117 545
rect 65 493 73 527
rect 107 493 117 527
rect 65 459 117 493
rect 65 425 73 459
rect 107 425 117 459
rect 65 391 117 425
rect 65 357 73 391
rect 107 357 117 391
rect 65 345 117 357
rect 147 533 201 545
rect 147 499 157 533
rect 191 499 201 533
rect 147 465 201 499
rect 147 431 157 465
rect 191 431 201 465
rect 147 345 201 431
rect 231 527 285 545
rect 231 493 241 527
rect 275 493 285 527
rect 231 459 285 493
rect 231 425 241 459
rect 275 425 285 459
rect 231 391 285 425
rect 231 357 241 391
rect 275 357 285 391
rect 231 345 285 357
rect 315 533 369 545
rect 315 499 325 533
rect 359 499 369 533
rect 315 465 369 499
rect 315 431 325 465
rect 359 431 369 465
rect 315 345 369 431
rect 399 511 453 545
rect 399 477 409 511
rect 443 477 453 511
rect 399 416 453 477
rect 399 382 409 416
rect 443 382 453 416
rect 399 345 453 382
rect 483 533 537 545
rect 483 499 493 533
rect 527 499 537 533
rect 483 465 537 499
rect 483 431 493 465
rect 527 431 537 465
rect 483 345 537 431
rect 567 511 621 545
rect 567 477 577 511
rect 611 477 621 511
rect 567 416 621 477
rect 567 382 577 416
rect 611 382 621 416
rect 567 345 621 382
rect 651 533 705 545
rect 651 499 661 533
rect 695 499 705 533
rect 651 465 705 499
rect 651 431 661 465
rect 695 431 705 465
rect 651 345 705 431
rect 735 511 789 545
rect 735 477 745 511
rect 779 477 789 511
rect 735 416 789 477
rect 735 382 745 416
rect 779 382 789 416
rect 735 345 789 382
rect 819 533 873 545
rect 819 499 829 533
rect 863 499 873 533
rect 819 465 873 499
rect 819 431 829 465
rect 863 431 873 465
rect 819 345 873 431
rect 903 511 957 545
rect 903 477 913 511
rect 947 477 957 511
rect 903 416 957 477
rect 903 382 913 416
rect 947 382 957 416
rect 903 345 957 382
rect 987 533 1039 545
rect 987 499 997 533
rect 1031 499 1039 533
rect 987 465 1039 499
rect 987 431 997 465
rect 1031 431 1039 465
rect 987 397 1039 431
rect 987 363 997 397
rect 1031 363 1039 397
rect 987 345 1039 363
<< ndiffc >>
rect 73 143 107 177
rect 157 111 191 145
rect 241 143 275 177
rect 325 111 359 145
rect 409 143 443 177
rect 493 111 527 145
rect 577 143 611 177
rect 661 111 695 145
rect 745 143 779 177
rect 829 111 863 145
rect 913 143 947 177
rect 997 175 1031 209
rect 997 107 1031 141
<< pdiffc >>
rect 73 493 107 527
rect 73 425 107 459
rect 73 357 107 391
rect 157 499 191 533
rect 157 431 191 465
rect 241 493 275 527
rect 241 425 275 459
rect 241 357 275 391
rect 325 499 359 533
rect 325 431 359 465
rect 409 477 443 511
rect 409 382 443 416
rect 493 499 527 533
rect 493 431 527 465
rect 577 477 611 511
rect 577 382 611 416
rect 661 499 695 533
rect 661 431 695 465
rect 745 477 779 511
rect 745 382 779 416
rect 829 499 863 533
rect 829 431 863 465
rect 913 477 947 511
rect 913 382 947 416
rect 997 499 1031 533
rect 997 431 1031 465
rect 997 363 1031 397
<< poly >>
rect 117 545 147 571
rect 201 545 231 571
rect 285 545 315 571
rect 369 545 399 571
rect 453 545 483 571
rect 537 545 567 571
rect 621 545 651 571
rect 705 545 735 571
rect 789 545 819 571
rect 873 545 903 571
rect 957 545 987 571
rect 117 309 147 345
rect 66 307 147 309
rect 201 307 231 345
rect 285 307 315 345
rect 66 297 315 307
rect 66 263 82 297
rect 116 263 150 297
rect 184 263 218 297
rect 252 263 315 297
rect 66 253 315 263
rect 66 251 147 253
rect 117 225 147 251
rect 201 225 231 253
rect 285 225 315 253
rect 369 307 399 345
rect 453 307 483 345
rect 537 307 567 345
rect 621 307 651 345
rect 705 307 735 345
rect 789 307 819 345
rect 873 307 903 345
rect 957 307 987 345
rect 369 297 987 307
rect 369 263 389 297
rect 423 263 457 297
rect 491 263 525 297
rect 559 263 593 297
rect 627 263 661 297
rect 695 263 729 297
rect 763 263 797 297
rect 831 263 987 297
rect 369 253 987 263
rect 369 225 399 253
rect 453 225 483 253
rect 537 225 567 253
rect 621 225 651 253
rect 705 225 735 253
rect 789 225 819 253
rect 873 225 903 253
rect 957 225 987 253
rect 117 69 147 95
rect 201 69 231 95
rect 285 69 315 95
rect 369 69 399 95
rect 453 69 483 95
rect 537 69 567 95
rect 621 69 651 95
rect 705 69 735 95
rect 789 69 819 95
rect 873 69 903 95
rect 957 69 987 95
<< polycont >>
rect 82 263 116 297
rect 150 263 184 297
rect 218 263 252 297
rect 389 263 423 297
rect 457 263 491 297
rect 525 263 559 297
rect 593 263 627 297
rect 661 263 695 297
rect 729 263 763 297
rect 797 263 831 297
<< locali >>
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 343 609
rect 377 575 435 609
rect 469 575 527 609
rect 561 575 619 609
rect 653 575 711 609
rect 745 575 803 609
rect 837 575 895 609
rect 929 575 987 609
rect 1021 575 1079 609
rect 1113 575 1142 609
rect 57 527 123 541
rect 57 493 73 527
rect 107 493 123 527
rect 57 459 123 493
rect 57 425 73 459
rect 107 425 123 459
rect 57 391 123 425
rect 157 533 191 575
rect 157 465 191 499
rect 157 415 191 431
rect 225 527 291 541
rect 225 493 241 527
rect 275 493 291 527
rect 225 459 291 493
rect 225 425 241 459
rect 275 425 291 459
rect 57 357 73 391
rect 107 371 123 391
rect 225 391 291 425
rect 325 533 359 575
rect 325 465 359 499
rect 325 415 359 431
rect 409 511 443 541
rect 409 416 443 477
rect 225 371 241 391
rect 107 357 241 371
rect 275 371 291 391
rect 477 533 543 575
rect 477 499 493 533
rect 527 499 543 533
rect 477 465 543 499
rect 477 431 493 465
rect 527 431 543 465
rect 477 415 543 431
rect 577 511 611 541
rect 577 416 611 477
rect 409 371 443 382
rect 645 533 711 575
rect 645 499 661 533
rect 695 499 711 533
rect 645 465 711 499
rect 645 431 661 465
rect 695 431 711 465
rect 645 415 711 431
rect 745 511 779 541
rect 745 416 779 477
rect 577 371 611 382
rect 813 533 879 575
rect 813 499 829 533
rect 863 499 879 533
rect 813 465 879 499
rect 813 431 829 465
rect 863 431 879 465
rect 813 415 879 431
rect 913 511 947 541
rect 913 416 947 477
rect 745 371 779 382
rect 913 371 947 382
rect 275 357 357 371
rect 57 337 357 357
rect 409 337 947 371
rect 981 533 1047 575
rect 981 499 997 533
rect 1031 499 1047 533
rect 981 465 1047 499
rect 981 431 997 465
rect 1031 431 1047 465
rect 981 397 1047 431
rect 981 363 997 397
rect 1031 363 1047 397
rect 981 345 1047 363
rect 66 297 286 303
rect 66 263 82 297
rect 116 263 150 297
rect 184 263 218 297
rect 252 263 286 297
rect 322 297 357 337
rect 322 263 389 297
rect 423 263 457 297
rect 491 263 525 297
rect 559 263 593 297
rect 627 263 661 297
rect 695 263 729 297
rect 763 263 797 297
rect 831 263 847 297
rect 322 229 357 263
rect 896 229 947 337
rect 73 195 357 229
rect 409 195 947 229
rect 73 177 107 195
rect 241 177 275 195
rect 73 99 107 143
rect 141 145 207 161
rect 141 111 157 145
rect 191 111 207 145
rect 141 65 207 111
rect 409 177 443 195
rect 241 100 275 143
rect 309 145 375 161
rect 309 111 325 145
rect 359 111 375 145
rect 309 65 375 111
rect 577 177 611 195
rect 409 99 443 143
rect 477 145 543 161
rect 477 111 493 145
rect 527 111 543 145
rect 477 65 543 111
rect 745 177 779 195
rect 577 99 611 143
rect 645 145 711 161
rect 645 111 661 145
rect 695 111 711 145
rect 645 65 711 111
rect 913 177 947 195
rect 745 99 779 143
rect 813 145 879 161
rect 813 111 829 145
rect 863 111 879 145
rect 813 65 879 111
rect 913 99 947 143
rect 981 209 1047 225
rect 981 175 997 209
rect 1031 175 1047 209
rect 981 141 1047 175
rect 981 107 997 141
rect 1031 107 1047 141
rect 981 65 1047 107
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 343 65
rect 377 31 435 65
rect 469 31 527 65
rect 561 31 619 65
rect 653 31 711 65
rect 745 31 803 65
rect 837 31 895 65
rect 929 31 987 65
rect 1021 31 1079 65
rect 1113 31 1142 65
<< viali >>
rect 67 575 101 609
rect 159 575 193 609
rect 251 575 285 609
rect 343 575 377 609
rect 435 575 469 609
rect 527 575 561 609
rect 619 575 653 609
rect 711 575 745 609
rect 803 575 837 609
rect 895 575 929 609
rect 987 575 1021 609
rect 1079 575 1113 609
rect 67 31 101 65
rect 159 31 193 65
rect 251 31 285 65
rect 343 31 377 65
rect 435 31 469 65
rect 527 31 561 65
rect 619 31 653 65
rect 711 31 745 65
rect 803 31 837 65
rect 895 31 929 65
rect 987 31 1021 65
rect 1079 31 1113 65
<< metal1 >>
rect 38 609 1142 640
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 343 609
rect 377 575 435 609
rect 469 575 527 609
rect 561 575 619 609
rect 653 575 711 609
rect 745 575 803 609
rect 837 575 895 609
rect 929 575 987 609
rect 1021 575 1079 609
rect 1113 575 1142 609
rect 38 544 1142 575
rect 38 65 1142 96
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 343 65
rect 377 31 435 65
rect 469 31 527 65
rect 561 31 619 65
rect 653 31 711 65
rect 745 31 803 65
rect 837 31 895 65
rect 929 31 987 65
rect 1021 31 1079 65
rect 1113 31 1142 65
rect 38 0 1142 31
<< labels >>
flabel locali s 252 269 286 303 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel locali s 896 201 930 235 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 896 269 930 303 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 160 269 194 303 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel locali s 68 31 102 65 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel locali s 68 575 102 609 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel locali s 896 337 930 371 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 68 269 102 303 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel pwell s 68 31 102 65 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 68 575 102 609 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 68 31 102 65 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 68 575 102 609 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 38 48 38 48 4 buf_8
<< properties >>
string FIXED_BBOX 38 48 1142 592
string path 0.190 0.240 5.710 0.240 
<< end >>
