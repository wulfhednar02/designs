magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -125 -200 1374 1540
<< l66d20 >>
rect 300 -200 500 1200
rect 265 1200 535 1530
<< l94d20 >>
rect 800 -125 1374 1125
<< l66d44 >>
rect 65 235 235 405
rect 65 595 235 765
rect 565 235 735 405
rect 565 595 735 765
rect 315 1280 485 1450
rect 940 235 1110 405
rect 940 595 1110 765
<< l67d44 >>
rect 65 235 235 405
rect 65 595 235 765
rect 565 235 735 405
rect 565 595 735 765
rect 315 1280 485 1450
<< l95d20 >>
rect 255 1190 545 1540
<< l67d20 >>
rect 65 155 235 845
rect 565 155 735 845
rect 235 1280 565 1450
rect 940 155 1110 845
<< l68d20 >>
rect 35 175 265 825
rect 535 175 765 825
rect 217 1250 583 1480
<< l65d20 >>
rect 0 0 800 1000
<< l93d44 >>
rect -125 -125 799 1125
<< l65d44 >>
rect 800 0 1250 1000
<< end >>
