magic
tech sky130A
magscale 1 2
timestamp 1699066547
<< pwell >>
rect -1 14 301 266
<< nmos >>
rect 85 40 125 240
<< ndiff >>
rect 25 193 85 240
rect 25 159 38 193
rect 72 159 85 193
rect 25 121 85 159
rect 25 87 38 121
rect 72 87 85 121
rect 25 40 85 87
rect 125 193 185 240
rect 125 159 138 193
rect 172 159 185 193
rect 125 121 185 159
rect 125 87 138 121
rect 172 87 185 121
rect 125 40 185 87
<< ndiffc >>
rect 38 159 72 193
rect 38 87 72 121
rect 138 159 172 193
rect 138 87 172 121
<< psubdiff >>
rect 185 193 275 240
rect 185 159 213 193
rect 247 159 275 193
rect 185 121 275 159
rect 185 87 213 121
rect 247 87 275 121
rect 185 40 275 87
<< psubdiffcont >>
rect 213 159 247 193
rect 213 87 247 121
<< poly >>
rect 78 330 132 346
rect 78 296 88 330
rect 122 296 132 330
rect 78 280 132 296
rect 85 240 125 280
rect 85 0 125 40
<< polycont >>
rect 88 296 122 330
<< locali >>
rect 72 296 88 330
rect 122 296 138 330
rect 38 193 72 209
rect 38 121 72 159
rect 38 71 72 87
rect 138 193 172 209
rect 138 121 172 159
rect 138 71 172 87
rect 213 193 247 209
rect 213 121 247 159
rect 213 71 247 87
<< viali >>
rect 88 296 122 330
rect 38 159 72 193
rect 38 87 72 121
rect 138 159 172 193
rect 138 87 172 121
<< metal1 >>
rect 68 330 142 336
rect 68 296 88 330
rect 122 296 142 330
rect 68 290 142 296
rect 32 193 78 205
rect 32 159 38 193
rect 72 159 78 193
rect 32 121 78 159
rect 32 87 38 121
rect 72 87 78 121
rect 32 75 78 87
rect 132 193 178 205
rect 132 159 138 193
rect 172 159 178 193
rect 132 121 178 159
rect 132 87 138 121
rect 172 87 178 121
rect 132 75 178 87
<< end >>
