magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -190 -240 1570 2960
<< l66d20 >>
rect 835 105 985 1060
rect 725 1060 995 1390
rect 835 1390 985 2615
rect 395 105 545 830
rect 365 830 545 950
rect 365 950 515 995
rect 135 995 515 1325
rect 365 1325 515 1500
rect 365 1500 545 1620
rect 395 1620 545 2615
<< l94d20 >>
rect 0 1420 1380 2910
<< l66d44 >>
rect 1035 445 1205 615
rect 1035 1810 1205 1980
rect 1035 2215 1205 2385
rect 775 1140 945 1310
rect 605 295 775 465
rect 605 1875 775 2045
rect 605 2215 775 2385
rect 185 1075 355 1245
rect 175 360 345 530
rect 175 1875 345 2045
rect 175 2215 345 2385
<< l67d44 >>
rect 1065 -85 1235 85
rect 1065 2635 1235 2805
rect 605 -85 775 85
rect 605 2635 775 2805
rect 145 -85 315 85
rect 145 2635 315 2805
<< l95d20 >>
rect 0 975 1380 1410
<< l67d20 >>
rect 1035 255 1295 760
rect 1115 760 1295 1560
rect 1025 1560 1295 2465
rect 0 -85 1380 85
rect 525 85 855 465
rect 175 255 345 635
rect 175 635 840 805
rect 670 805 840 1060
rect 670 1060 945 1390
rect 670 1390 840 1535
rect 165 1535 840 1705
rect 165 1705 345 2465
rect 525 1875 855 2635
rect 0 2635 1380 2805
rect 105 985 445 1355
<< l68d20 >>
rect 0 -240 1380 240
rect 0 2480 1380 2960
<< l65d20 >>
rect 135 235 1245 755
rect 135 1695 1245 2485
<< l93d44 >>
rect 0 -190 1380 1015
<< l64d20 >>
rect -190 1305 1570 2910
<< l68d16 >>
rect 155 -85 325 85
rect 145 2635 315 2805
<< l236d0 >>
rect 0 0 1380 2720
<< l122d16 >>
rect 155 -85 325 85
<< l64d16 >>
rect 145 2635 315 2805
<< l81d4 >>
rect 0 0 1380 2720
<< l78d44 >>
rect 0 1250 1380 2720
<< l67d16 >>
rect 1055 425 1225 595
rect 1055 1785 1225 1955
rect 1055 2125 1225 2295
rect 145 1105 315 1275
rect 145 2635 315 2805
rect 155 -85 325 85
<< labels >>
rlabel l67d5 230 2720 230 2720 0 VPWR
rlabel l67d5 230 0 230 0 0 VGND
rlabel l67d5 1140 510 1140 510 0 X
rlabel l67d5 1140 1870 1140 1870 0 X
rlabel l67d5 1140 2210 1140 2210 0 X
rlabel l67d5 230 1190 230 1190 0 A
rlabel l64d59 230 0 230 0 0 VNB
rlabel l64d5 230 2720 230 2720 0 VPB
rlabel l68d5 230 0 230 0 0 VGND
rlabel l68d5 230 2720 230 2720 0 VPWR
rlabel l83d44 0 0 0 0 0 buf_1
<< end >>
