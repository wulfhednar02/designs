magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -190 -240 5710 2960
<< l66d20 >>
rect 395 105 545 1015
rect 140 1015 545 1025
rect 815 105 965 1025
rect 1235 105 1385 1025
rect 140 1025 1385 1295
rect 140 1295 545 1305
rect 395 1305 545 2615
rect 815 1295 965 2615
rect 1235 1295 1385 2615
rect 1655 105 1805 1025
rect 2075 105 2225 1025
rect 2495 105 2645 1025
rect 2915 105 3065 1025
rect 3335 105 3485 1025
rect 3755 105 3905 1025
rect 4175 105 4325 1025
rect 4595 105 4745 1025
rect 1655 1025 4745 1295
rect 1655 1295 1805 2615
rect 2075 1295 2225 2615
rect 2495 1295 2645 2615
rect 2915 1295 3065 2615
rect 3335 1295 3485 2615
rect 3755 1295 3905 2615
rect 4175 1295 4325 2615
rect 4595 1295 4745 2615
<< l94d20 >>
rect 0 1355 5520 2910
<< l66d44 >>
rect 4795 1575 4965 1745
rect 4795 635 4965 805
rect 4795 295 4965 465
rect 3115 315 3285 485
rect 3455 1075 3625 1245
rect 3535 1670 3705 1840
rect 3535 475 3705 645
rect 3115 1915 3285 2085
rect 2695 1670 2865 1840
rect 2275 1915 2445 2085
rect 4795 1915 4965 2085
rect 3955 2255 4125 2425
rect 3955 1915 4125 2085
rect 3955 315 4125 485
rect 4375 2145 4545 2315
rect 4375 1670 4545 1840
rect 175 2225 345 2395
rect 175 1885 345 2055
rect 175 1545 345 1715
rect 175 475 345 645
rect 220 1075 390 1245
rect 560 1075 730 1245
rect 595 2255 765 2425
rect 595 1915 765 2085
rect 595 315 765 485
rect 900 1075 1070 1245
rect 1015 2225 1185 2395
rect 1015 1885 1185 2055
rect 1015 1545 1185 1715
rect 1015 475 1185 645
rect 1435 2255 1605 2425
rect 1435 1915 1605 2085
rect 1435 315 1605 485
rect 1755 1075 1925 1245
rect 1855 2145 2025 2315
rect 1855 1670 2025 1840
rect 4375 475 4545 645
rect 4795 2255 4965 2425
rect 1855 475 2025 645
rect 2095 1075 2265 1245
rect 2275 2255 2445 2425
rect 2275 315 2445 485
rect 2435 1075 2605 1245
rect 2695 2145 2865 2315
rect 2695 475 2865 645
rect 2775 1075 2945 1245
rect 3115 2255 3285 2425
rect 3115 1075 3285 1245
rect 3795 1075 3965 1245
rect 3535 2145 3705 2315
<< l67d44 >>
rect 145 2635 315 2805
rect 145 -85 315 85
rect 605 2635 775 2805
rect 605 -85 775 85
rect 1065 2635 1235 2805
rect 1065 -85 1235 85
rect 1525 2635 1695 2805
rect 1525 -85 1695 85
rect 1985 2635 2155 2805
rect 1985 -85 2155 85
rect 2445 2635 2615 2805
rect 2445 -85 2615 85
rect 2905 2635 3075 2805
rect 2905 -85 3075 85
rect 3365 2635 3535 2805
rect 3365 -85 3535 85
rect 3825 2635 3995 2805
rect 3825 -85 3995 85
rect 4285 2635 4455 2805
rect 4285 -85 4455 85
rect 4745 2635 4915 2805
rect 4745 -85 4915 85
rect 5205 2635 5375 2805
rect 5205 -85 5375 85
<< l95d20 >>
rect 0 975 5520 1345
<< l67d20 >>
rect 175 255 345 735
rect 1015 260 1185 735
rect 175 735 1595 905
rect 1420 905 1595 1075
rect 1420 1075 4045 1245
rect 1420 1245 1595 1445
rect 95 1445 1595 1615
rect 95 1615 425 2465
rect 935 1615 1265 2465
rect 0 -85 5520 85
rect 515 85 845 565
rect 1355 85 1685 565
rect 2195 85 2525 565
rect 3035 85 3365 565
rect 3875 85 4205 565
rect 4715 85 5045 885
rect 595 1835 765 2635
rect 1435 1835 1605 2635
rect 2195 1835 2525 2635
rect 3035 1835 3365 2635
rect 3875 1835 4205 2635
rect 4715 1485 5045 2635
rect 0 2635 5520 2805
rect 1855 255 2025 735
rect 2695 255 2865 735
rect 3535 255 3705 735
rect 4375 255 4545 735
rect 1855 735 4545 905
rect 4290 905 4545 1445
rect 1855 1445 4545 1615
rect 1855 1615 2025 2465
rect 2695 1615 2865 2465
rect 3535 1615 3705 2465
rect 4375 1615 4545 2465
rect 140 1075 1240 1275
<< l68d20 >>
rect 0 2480 5520 2960
rect 0 -240 5520 240
<< l65d20 >>
rect 135 1485 5005 2485
rect 135 235 5005 885
<< l93d44 >>
rect 0 -190 5520 1015
<< l64d20 >>
rect -190 1305 5710 2910
<< l68d16 >>
rect 150 -85 320 85
rect 150 2635 320 2805
<< l236d0 >>
rect 0 0 5520 2720
<< l122d16 >>
rect 150 -85 320 85
<< l64d16 >>
rect 150 2635 320 2805
<< l81d4 >>
rect 0 0 5520 2720
<< l78d44 >>
rect 0 1250 5520 2720
<< l67d16 >>
rect 150 1105 320 1275
rect 610 1105 780 1275
rect 1070 1105 1240 1275
rect 4290 1445 4460 1615
rect 4290 1105 4460 1275
rect 4290 765 4460 935
rect 150 -85 320 85
rect 150 2635 320 2805
<< labels >>
rlabel l67d5 1155 1190 1155 1190 0 A
rlabel l67d5 4375 850 4375 850 0 X
rlabel l67d5 4375 1190 4375 1190 0 X
rlabel l67d5 695 1190 695 1190 0 A
rlabel l67d5 230 0 230 0 0 VGND
rlabel l67d5 235 2720 235 2720 0 VPWR
rlabel l67d5 4375 1530 4375 1530 0 X
rlabel l67d5 235 1190 235 1190 0 A
rlabel l64d59 235 0 235 0 0 VNB
rlabel l64d5 235 2720 235 2720 0 VPB
rlabel l68d5 230 0 230 0 0 VGND
rlabel l68d5 235 2720 235 2720 0 VPWR
rlabel l83d44 0 0 0 0 0 buf_8
<< end >>
