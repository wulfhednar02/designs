magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< error_s >>
rect 968 4527 1037 4596
rect 1038 4527 1108 4554
rect 1109 4527 1178 4596
rect 968 4526 1178 4527
rect 606 4525 784 4526
rect 854 4525 1107 4526
rect 1108 4525 1540 4526
rect 606 4484 784 4485
rect 854 4484 1037 4485
rect 1038 4484 1107 4485
rect 1109 4484 1540 4485
rect 1222 4030 1291 4099
rect 1292 4030 1362 4057
rect 1363 4030 1432 4099
rect 1222 4029 1432 4030
rect 860 4028 1361 4029
rect 1362 4028 1794 4029
rect 860 3987 1291 3988
rect 1292 3987 1361 3988
rect 1363 3987 1794 3988
rect 968 3533 1037 3602
rect 1038 3533 1108 3560
rect 1109 3533 1178 3602
rect 968 3532 1178 3533
rect 606 3531 1107 3532
rect 1108 3531 1540 3532
rect 606 3490 1037 3491
rect 1038 3490 1107 3491
rect 1109 3490 1540 3491
rect 1222 3036 1291 3105
rect 1292 3036 1362 3063
rect 1363 3036 1432 3105
rect 1222 3035 1432 3036
rect 860 3034 1361 3035
rect 1362 3034 1794 3035
rect 860 2993 1291 2994
rect 1292 2993 1361 2994
rect 1363 2993 1794 2994
rect 968 2539 1037 2608
rect 1038 2539 1108 2566
rect 1109 2539 1178 2608
rect 968 2538 1178 2539
rect 606 2537 1107 2538
rect 1108 2537 1540 2538
rect 606 2496 1037 2497
rect 1038 2496 1107 2497
rect 1109 2496 1540 2497
rect 1222 2042 1291 2111
rect 1292 2042 1362 2069
rect 1363 2042 1432 2111
rect 1222 2041 1432 2042
rect 860 2040 1361 2041
rect 1362 2040 1794 2041
rect 860 1999 1291 2000
rect 1292 1999 1361 2000
rect 1363 1999 1794 2000
rect 968 1545 1037 1614
rect 1038 1545 1108 1572
rect 1109 1545 1178 1614
rect 968 1544 1178 1545
rect 606 1543 1107 1544
rect 1108 1543 1540 1544
rect 606 1502 1037 1503
rect 1038 1502 1107 1503
rect 1109 1502 1540 1503
rect 1222 1048 1291 1117
rect 1292 1048 1362 1075
rect 1363 1048 1432 1117
rect 1222 1047 1432 1048
rect 860 1046 1361 1047
rect 1362 1046 1794 1047
rect 860 1005 1291 1006
rect 1292 1005 1361 1006
rect 1363 1005 1794 1006
<< metal1 >>
rect 794 4585 844 5006
rect 1041 4952 1105 4958
rect 1041 4900 1047 4952
rect 1099 4900 1105 4952
rect 1041 4880 1105 4900
rect 1041 4828 1047 4880
rect 1099 4828 1105 4880
rect 1041 4808 1105 4828
rect 1041 4756 1047 4808
rect 1099 4756 1105 4808
rect 1041 4736 1105 4756
rect 1041 4684 1047 4736
rect 1099 4684 1105 4736
rect 1041 4664 1105 4684
rect 1041 4612 1047 4664
rect 1099 4612 1105 4664
rect 1041 4592 1105 4612
rect 1041 4540 1047 4592
rect 1099 4540 1105 4592
rect 1041 4534 1105 4540
rect 540 4088 590 4509
rect 794 4038 1352 4475
rect 286 3591 336 4012
rect 540 3541 1352 3978
rect 32 3094 82 3515
rect 286 3044 1352 3481
rect 32 2547 1352 2984
rect 32 2050 1352 2487
rect 32 1519 82 1940
rect 286 1553 1352 1990
rect 286 1022 336 1443
rect 540 1056 1352 1493
rect 540 525 590 946
rect 794 559 1352 996
rect 794 28 844 449
rect 1041 445 1105 451
rect 1041 393 1047 445
rect 1099 393 1105 445
rect 1041 373 1105 393
rect 1041 321 1047 373
rect 1099 321 1105 373
rect 1041 301 1105 321
rect 1041 249 1047 301
rect 1099 249 1105 301
rect 1041 229 1105 249
rect 1041 177 1047 229
rect 1099 177 1105 229
rect 1041 157 1105 177
rect 1041 105 1047 157
rect 1099 105 1105 157
rect 1041 85 1105 105
rect 1041 33 1047 85
rect 1099 33 1105 85
rect 1041 27 1105 33
<< via1 >>
rect 1047 4900 1099 4952
rect 1047 4828 1099 4880
rect 1047 4756 1099 4808
rect 1047 4684 1099 4736
rect 1047 4612 1099 4664
rect 1047 4540 1099 4592
rect 1047 393 1099 445
rect 1047 321 1099 373
rect 1047 249 1099 301
rect 1047 177 1099 229
rect 1047 105 1099 157
rect 1047 33 1099 85
<< metal2 >>
rect 1041 4952 1105 4958
rect 1041 4900 1047 4952
rect 1099 4900 1105 4952
rect 1041 4880 1105 4900
rect 1041 4828 1047 4880
rect 1099 4828 1105 4880
rect 1041 4808 1105 4828
rect 1041 4756 1047 4808
rect 1099 4756 1105 4808
rect 1041 4736 1105 4756
rect 1041 4684 1047 4736
rect 1099 4684 1105 4736
rect 1041 4664 1105 4684
rect 1041 4612 1047 4664
rect 1099 4612 1105 4664
rect 1041 4592 1105 4612
rect 1041 4540 1047 4592
rect 1099 4540 1105 4592
rect 1041 4534 1105 4540
rect 1041 445 1105 451
rect 1041 393 1047 445
rect 1099 393 1105 445
rect 1041 373 1105 393
rect 1041 321 1047 373
rect 1099 321 1105 373
rect 1041 301 1105 321
rect 1041 249 1047 301
rect 1099 249 1105 301
rect 1041 229 1105 249
rect 1041 177 1047 229
rect 1099 177 1105 229
rect 1041 157 1105 177
rect 1041 105 1047 157
rect 1099 105 1105 157
rect 1041 85 1105 105
rect 1041 33 1047 85
rect 1099 33 1105 85
rect 1041 27 1105 33
use res_poly$3  res_poly$3_0
timestamp 1698900908
transform 1 0 565 0 1 1001
box -35 -482 35 482
use res_poly$3  res_poly$3_1
timestamp 1698900908
transform 1 0 819 0 1 504
box -35 -482 35 482
use res_poly$3  res_poly$3_2
timestamp 1698900908
transform 1 0 565 0 1 4033
box -35 -482 35 482
use res_poly$3  res_poly$3_3
timestamp 1698900908
transform 1 0 819 0 1 4530
box -35 -482 35 482
use res_poly$3  res_poly$3_4
timestamp 1698900908
transform 1 0 1073 0 1 504
box -35 -482 35 482
use res_poly$3  res_poly$3_5
timestamp 1698900908
transform 1 0 57 0 1 1995
box -35 -482 35 482
use res_poly$3  res_poly$3_6
timestamp 1698900908
transform 1 0 311 0 1 3536
box -35 -482 35 482
use res_poly$3  res_poly$3_7
timestamp 1698900908
transform 1 0 311 0 1 1498
box -35 -482 35 482
use res_poly$3  res_poly$3_8
timestamp 1698900908
transform 1 0 57 0 1 3039
box -35 -482 35 482
use res_poly$4  res_poly$4_0
timestamp 1698900908
transform 1 0 1327 0 1 2020
box -467 -458 467 458
use res_poly$4  res_poly$4_1
timestamp 1698900908
transform 1 0 1073 0 1 4505
box -467 -458 467 458
use res_poly$4  res_poly$4_2
timestamp 1698900908
transform 1 0 1073 0 1 3511
box -467 -458 467 458
use res_poly$4  res_poly$4_3
timestamp 1698900908
transform 1 0 1327 0 1 4008
box -467 -458 467 458
use res_poly$4  res_poly$4_4
timestamp 1698900908
transform 1 0 1327 0 1 3014
box -467 -458 467 458
use res_poly$4  res_poly$4_5
timestamp 1698900908
transform 1 0 1327 0 1 1026
box -467 -458 467 458
use res_poly$4  res_poly$4_6
timestamp 1698900908
transform 1 0 1073 0 1 1523
box -467 -458 467 458
use res_poly$4  res_poly$4_7
timestamp 1698900908
transform 1 0 1073 0 1 2517
box -467 -458 467 458
<< labels >>
flabel metal1 s 794 4038 1352 4474 0 FreeSans 44 0 0 0 OUT
port 2 nsew
flabel metal1 s 937 4260 937 4260 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 923 4449 923 4449 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 286 3591 336 4012 0 FreeSans 44 0 0 0 DAC5
port 3 nsew
flabel metal1 s 311 3804 311 3804 0 FreeSans 44 0 0 0 DAC5
flabel metal1 s 308 3984 308 3984 0 FreeSans 44 0 0 0 DAC5
flabel metal1 s 540 4088 590 4509 0 FreeSans 44 0 0 0 DAC6
port 4 nsew
flabel metal1 s 794 4585 844 5006 0 FreeSans 44 0 0 0 DAC7
port 5 nsew
flabel metal1 s 563 4481 563 4481 0 FreeSans 44 0 0 0 DAC6
flabel metal1 s 565 4296 565 4296 0 FreeSans 44 0 0 0 DAC6
flabel metal1 s 817 4615 817 4615 0 FreeSans 44 0 0 0 DAC7
flabel metal1 s 817 4796 817 4796 0 FreeSans 44 0 0 0 DAC7
flabel metal1 s 1196 4438 1196 4438 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 1195 4273 1195 4273 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 1196 4080 1196 4080 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 32 3094 82 3515 0 FreeSans 44 0 0 0 DAC4
port 6 nsew
flabel metal1 s 55 3304 55 3304 0 FreeSans 44 0 0 0 DAC4
flabel metal1 s 55 3124 55 3124 0 FreeSans 44 0 0 0 DAC4
flabel metal1 s 32 1519 82 1939 0 FreeSans 44 0 0 0 DAC3
port 7 nsew
flabel metal1 s 58 1735 58 1735 0 FreeSans 44 0 0 0 DAC3
flabel metal1 s 56 1550 56 1550 0 FreeSans 44 0 0 0 DAC3
flabel metal1 s 286 1022 336 1442 0 FreeSans 44 0 0 0 DAC2
port 8 nsew
flabel metal1 s 309 1411 309 1411 0 FreeSans 44 0 0 0 DAC2
flabel metal1 s 312 1054 312 1054 0 FreeSans 44 0 0 0 DAC2
flabel metal1 s 540 525 590 945 0 FreeSans 44 0 0 0 DAC1
port 9 nsew
flabel metal1 s 568 919 568 919 0 FreeSans 44 0 0 0 DAC1
flabel metal1 s 566 556 566 556 0 FreeSans 44 0 0 0 DAC1
flabel metal1 s 794 28 844 448 0 FreeSans 44 0 0 0 DAC0
port 10 nsew
flabel metal1 s 818 419 818 419 0 FreeSans 44 0 0 0 DAC0
flabel metal1 s 818 59 818 59 0 FreeSans 44 0 0 0 DAC0
flabel metal2 s 1041 4534 1105 4958 0 FreeSans 44 0 0 0 VDD
port 12 nsew
flabel metal2 s 1072 4749 1072 4749 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 1072 4565 1072 4565 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 1041 27 1105 451 0 FreeSans 44 0 0 0 VSS
port 13 nsew
flabel metal2 s 1070 57 1070 57 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 1071 418 1071 418 0 FreeSans 44 0 0 0 VSS
<< end >>
