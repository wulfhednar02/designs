magic
tech sky130A
timestamp 1698900908
<< end >>
