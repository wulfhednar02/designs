magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< error_s >>
rect 17141 21212 17153 21218
rect 17163 21194 17165 21206
rect 20416 21122 20422 21128
rect 20386 21098 20392 21118
rect 20344 21010 20350 21030
rect 20386 20988 20392 20994
rect 17163 20826 17165 20838
rect 17141 20814 17153 20820
rect 2298 20388 2498 20410
rect 21916 20398 21944 20468
rect 22910 20398 22938 20468
rect 23904 20398 23932 20468
rect 24898 20398 24926 20468
rect 22413 20144 22441 20214
rect 23407 20144 23435 20214
rect 24401 20144 24429 20214
rect 25395 20144 25423 20214
rect 11340 20008 11540 20030
rect 2288 19666 8340 19667
rect 11330 19286 17382 19287
rect 21302 17852 21345 17920
rect 1317 9586 1339 9824
rect 2006 9586 2049 15654
rect 21344 11826 21345 17852
rect 22066 17668 22088 17868
rect 2006 9560 2007 9586
rect 2527 1366 2549 1604
rect 3216 1366 3259 7434
rect 14969 4073 21105 4116
rect 4668 3749 4811 4003
rect 4922 2154 5065 3749
rect 20799 3384 21037 3406
rect 6930 2154 13066 2197
rect 12760 1465 12998 1487
rect 3216 1340 3217 1366
<< metal1 >>
rect 1856 20837 11335 21274
rect 400 20400 2293 20837
rect 400 9565 836 20400
rect 1856 17575 2264 20197
rect 10898 20020 11335 20837
rect 16983 21212 17057 21786
rect 21755 21726 22025 21786
rect 22252 21726 22577 21786
rect 22749 21726 23129 21786
rect 23246 21726 23681 21786
rect 24159 21726 24521 21786
rect 24711 21726 25018 21786
rect 25263 21726 25514 21786
rect 25815 21726 26012 21786
rect 16983 20820 17108 21212
rect 20526 21018 20645 21092
rect 10303 19409 11191 19817
rect 20571 19437 20645 21018
rect 21755 20772 21815 21726
rect 22252 21026 22312 21726
rect 22749 21280 22809 21726
rect 23246 21534 23306 21726
rect 24461 21534 24521 21726
rect 22885 21474 23306 21534
rect 24460 21474 24881 21534
rect 24958 21280 25018 21726
rect 22388 21220 22809 21280
rect 24957 21220 25378 21280
rect 25455 21026 25515 21726
rect 21891 20966 22312 21026
rect 25454 20966 25875 21026
rect 25952 20772 26012 21726
rect 21394 20712 21815 20772
rect 25951 20712 26372 20772
rect 19345 19029 20645 19437
rect 20291 18017 20571 19029
rect 21926 18310 22362 20154
rect 21926 17873 22964 18310
rect 400 9128 1273 9565
rect 1476 9128 3474 9536
rect 836 1345 1273 9128
rect 836 908 2483 1345
rect 5009 1316 5417 2004
rect 13048 1624 13456 3923
rect 21087 3543 21495 9863
rect 22528 3340 22964 17873
rect 21058 2903 22964 3340
rect 21058 1421 21495 2903
rect 2686 1016 5417 1316
rect 13019 984 21495 1421
rect 13019 908 13456 984
rect 2046 472 13456 908
<< metal2 >>
rect 0 21370 3864 22304
rect 27916 22260 31464 22304
rect 8702 21370 16506 22084
rect 27916 21370 31116 22260
rect 0 21116 31116 21370
rect 0 20290 16692 21116
rect 20897 20828 31116 21116
rect 20897 20290 21026 20828
rect 21437 20462 21871 20470
rect 21437 20406 21446 20462
rect 21502 20406 21536 20462
rect 21592 20406 21626 20462
rect 21682 20406 21716 20462
rect 21772 20406 21806 20462
rect 21862 20406 21871 20462
rect 21437 20396 21871 20406
rect 0 20006 21026 20290
rect 22225 20006 31116 20828
rect 0 18754 31116 20006
rect 0 17854 1919 18754
rect 10697 18393 31116 18754
rect 0 9252 2904 17854
rect 10697 17755 10970 18393
rect 3909 17367 10970 17755
rect 3909 9770 19400 17367
rect 3909 9252 4122 9770
rect 5132 9462 19400 9770
rect 20449 9462 31116 18393
rect 0 1079 4122 9252
rect 5132 5988 31116 9462
rect 5132 4955 12636 5988
rect 21449 4956 31116 5988
rect 13400 4955 31116 4956
rect 5132 4086 31116 4955
rect 13400 3056 31116 4086
rect 5132 1079 31116 3056
rect 0 44 31116 1079
rect 31412 44 31464 22260
rect 0 0 31464 44
<< via2 >>
rect 17126 20716 17182 20772
rect 17206 20716 17262 20772
rect 17286 20716 17342 20772
rect 17366 20716 17422 20772
rect 17446 20716 17502 20772
rect 17526 20716 17582 20772
rect 17606 20716 17662 20772
rect 17686 20716 17742 20772
rect 17766 20716 17822 20772
rect 17846 20716 17902 20772
rect 17926 20716 17982 20772
rect 18006 20716 18062 20772
rect 18086 20716 18142 20772
rect 18166 20716 18222 20772
rect 18246 20716 18302 20772
rect 18326 20716 18382 20772
rect 18406 20716 18462 20772
rect 18486 20716 18542 20772
rect 18566 20716 18622 20772
rect 18646 20716 18702 20772
rect 18726 20716 18782 20772
rect 18806 20716 18862 20772
rect 18886 20716 18942 20772
rect 18966 20716 19022 20772
rect 19046 20716 19102 20772
rect 19126 20716 19182 20772
rect 19206 20716 19262 20772
rect 19286 20716 19342 20772
rect 19366 20716 19422 20772
rect 19446 20716 19502 20772
rect 19526 20716 19582 20772
rect 19606 20716 19662 20772
rect 19686 20716 19742 20772
rect 19766 20716 19822 20772
rect 19846 20716 19902 20772
rect 19926 20716 19982 20772
rect 20006 20716 20062 20772
rect 20086 20716 20142 20772
rect 20166 20716 20222 20772
rect 20246 20716 20302 20772
rect 20326 20716 20382 20772
rect 20406 20716 20462 20772
rect 21446 20406 21502 20462
rect 21536 20406 21592 20462
rect 21626 20406 21682 20462
rect 21716 20406 21772 20462
rect 21806 20406 21862 20462
rect 2366 18198 10262 18334
rect 11408 17818 19304 17954
rect 3340 9638 3476 17534
rect 19875 9904 20011 17800
rect 4550 1418 4686 9314
rect 13089 5406 20985 5542
rect 5050 3488 12946 3624
rect 31116 44 31412 22260
<< metal3 >>
rect 0 22264 8226 22304
rect 0 40 48 22264
rect 352 21370 8226 22264
rect 27916 21370 30633 22304
rect 352 20772 30633 21370
rect 352 20716 17126 20772
rect 17182 20716 17206 20772
rect 17262 20716 17286 20772
rect 17342 20716 17366 20772
rect 17422 20716 17446 20772
rect 17502 20716 17526 20772
rect 17582 20716 17606 20772
rect 17662 20716 17686 20772
rect 17742 20716 17766 20772
rect 17822 20716 17846 20772
rect 17902 20716 17926 20772
rect 17982 20716 18006 20772
rect 18062 20716 18086 20772
rect 18142 20716 18166 20772
rect 18222 20716 18246 20772
rect 18302 20716 18326 20772
rect 18382 20716 18406 20772
rect 18462 20716 18486 20772
rect 18542 20716 18566 20772
rect 18622 20716 18646 20772
rect 18702 20716 18726 20772
rect 18782 20716 18806 20772
rect 18862 20716 18886 20772
rect 18942 20716 18966 20772
rect 19022 20716 19046 20772
rect 19102 20716 19126 20772
rect 19182 20716 19206 20772
rect 19262 20716 19286 20772
rect 19342 20716 19366 20772
rect 19422 20716 19446 20772
rect 19502 20716 19526 20772
rect 19582 20716 19606 20772
rect 19662 20716 19686 20772
rect 19742 20716 19766 20772
rect 19822 20716 19846 20772
rect 19902 20716 19926 20772
rect 19982 20716 20006 20772
rect 20062 20716 20086 20772
rect 20142 20716 20166 20772
rect 20222 20716 20246 20772
rect 20302 20716 20326 20772
rect 20382 20716 20406 20772
rect 20462 20716 30633 20772
rect 352 20462 30633 20716
rect 352 20406 21446 20462
rect 21502 20406 21536 20462
rect 21592 20406 21626 20462
rect 21682 20406 21716 20462
rect 21772 20406 21806 20462
rect 21862 20406 30633 20462
rect 352 18334 30633 20406
rect 352 18198 2366 18334
rect 10262 18198 30633 18334
rect 352 17954 30633 18198
rect 352 17818 11408 17954
rect 19304 17818 30633 17954
rect 352 17800 30633 17818
rect 352 17534 19875 17800
rect 352 9638 3340 17534
rect 3476 9904 19875 17534
rect 20011 9904 30633 17800
rect 3476 9638 30633 9904
rect 352 9314 30633 9638
rect 352 1418 4550 9314
rect 4686 5542 30633 9314
rect 4686 5406 13089 5542
rect 20985 5406 30633 5542
rect 4686 3624 30633 5406
rect 4686 3488 5050 3624
rect 12946 3488 30633 3624
rect 4686 1418 30633 3488
rect 352 40 30633 1418
rect 0 0 30633 40
rect 31064 22264 31464 22304
rect 31064 40 31112 22264
rect 31416 40 31464 22264
rect 31064 0 31464 40
<< via3 >>
rect 48 40 352 22264
rect 31112 22260 31416 22264
rect 31112 44 31116 22260
rect 31116 44 31412 22260
rect 31412 44 31416 22260
rect 31112 40 31416 44
<< metal4 >>
rect 0 22264 400 22304
rect 0 40 48 22264
rect 352 40 400 22264
rect 4294 22104 4354 22304
rect 4846 22104 4906 22304
rect 5398 22104 5458 22304
rect 5950 22104 6010 22304
rect 6502 22104 6562 22304
rect 7054 22104 7114 22304
rect 7606 22104 7666 22304
rect 8158 22104 8218 22304
rect 8710 22104 8770 22304
rect 9262 22104 9322 22304
rect 9814 22104 9874 22304
rect 10366 22104 10426 22304
rect 10918 22104 10978 22304
rect 11470 22104 11530 22304
rect 12022 22104 12082 22304
rect 12574 22104 12634 22304
rect 13126 22104 13186 22304
rect 13678 22104 13738 22304
rect 14230 22104 14290 22304
rect 14782 22104 14842 22304
rect 15334 22104 15394 22304
rect 15886 22104 15946 22304
rect 16438 22104 16498 22304
rect 16990 22104 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22104 22018 22304
rect 22510 22104 22570 22304
rect 23062 22104 23122 22304
rect 23614 22104 23674 22304
rect 24166 22104 24226 22304
rect 24718 22104 24778 22304
rect 25270 22104 25330 22304
rect 25822 22104 25882 22304
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 31064 22264 31464 22304
rect 0 0 400 40
rect 31064 40 31112 22264
rect 31416 40 31464 22264
rect 31064 0 31464 40
use dac_8bit  dac_8bit_0
timestamp 1698982078
transform 0 -1 26418 -1 0 21576
box 92 40 1432 5030
use driver  driver_0
timestamp 1698982078
transform -1 0 20538 0 -1 21336
box 0 0 3485 640
use inv_strvd  inv_strvd_0
timestamp 1698982078
transform 0 1 2220 1 0 1201
box 0 -1 8241 2591
use inv_strvd  inv_strvd_1
timestamp 1698982078
transform 1 0 2149 0 -1 20663
box 0 -1 8241 2591
use inv_strvd  inv_strvd_2
timestamp 1698982078
transform 1 0 11191 0 -1 20283
box 0 -1 8241 2591
use inv_strvd  inv_strvd_3
timestamp 1698982078
transform -1 0 13163 0 1 1158
box 0 -1 8241 2591
use inv_strvd  inv_strvd_4
timestamp 1698982078
transform 0 -1 22341 -1 0 18017
box 0 -1 8241 2591
use inv_strvd  inv_strvd_5
timestamp 1698982078
transform 0 1 1010 1 0 9421
box 0 -1 8241 2591
use inv_strvd  inv_strvd_6
timestamp 1698982078
transform -1 0 21202 0 1 3077
box 0 -1 8241 2591
use pin_connect  pin_connect_0
timestamp 1698982078
transform 1 0 27470 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_1
timestamp 1698982078
transform 1 0 26918 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_2
timestamp 1698982078
transform 1 0 26366 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_3
timestamp 1698982078
transform 1 0 25814 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_4
timestamp 1698982078
transform 1 0 25262 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_5
timestamp 1698982078
transform 1 0 24710 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_6
timestamp 1698982078
transform 1 0 24158 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_7
timestamp 1698982078
transform 1 0 23606 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_8
timestamp 1698982078
transform 1 0 23054 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_9
timestamp 1698982078
transform 1 0 22502 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_10
timestamp 1698982078
transform 1 0 21950 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_11
timestamp 1698982078
transform 1 0 21398 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_12
timestamp 1698982078
transform 1 0 20846 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_13
timestamp 1698982078
transform 1 0 20294 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_14
timestamp 1698982078
transform 1 0 19742 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_15
timestamp 1698982078
transform 1 0 19190 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_16
timestamp 1698982078
transform 1 0 18638 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_17
timestamp 1698982078
transform 1 0 18086 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_18
timestamp 1698982078
transform 1 0 17534 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_19
timestamp 1698982078
transform 1 0 16982 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_20
timestamp 1698982078
transform 1 0 16430 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_21
timestamp 1698982078
transform 1 0 15878 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_22
timestamp 1698982078
transform 1 0 15326 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_23
timestamp 1698982078
transform 1 0 14774 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_24
timestamp 1698982078
transform 1 0 14222 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_25
timestamp 1698982078
transform 1 0 13670 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_26
timestamp 1698982078
transform 1 0 13118 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_27
timestamp 1698982078
transform 1 0 12566 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_28
timestamp 1698982078
transform 1 0 12014 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_29
timestamp 1698982078
transform 1 0 11462 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_30
timestamp 1698982078
transform 1 0 10910 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_31
timestamp 1698982078
transform 1 0 10358 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_32
timestamp 1698982078
transform 1 0 9806 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_33
timestamp 1698982078
transform 1 0 9254 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_34
timestamp 1698982078
transform 1 0 8702 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_35
timestamp 1698982078
transform 1 0 8150 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_36
timestamp 1698982078
transform 1 0 7598 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_37
timestamp 1698982078
transform 1 0 7046 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_38
timestamp 1698982078
transform 1 0 6494 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_39
timestamp 1698982078
transform 1 0 5942 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_40
timestamp 1698982078
transform 1 0 5390 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_41
timestamp 1698982078
transform 1 0 4838 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_42
timestamp 1698982078
transform 1 0 4286 0 1 21786
box 0 0 76 518
use tt_um_template  tt_um_template_0
timestamp 1698982078
transform 1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel metal4 s 31064 0 31464 22304 0 FreeSans 2000 0 0 0 VGND
port 2 nsew
rlabel metal4 s 26926 22104 26986 22304 4 clk
port 3 nsew
rlabel metal4 s 27478 22104 27538 22304 4 ena
port 4 nsew
rlabel metal4 s 26374 22104 26434 22304 4 rst_n
port 5 nsew
rlabel metal4 s 25822 22104 25882 22304 4 ui_in[0]
port 6 nsew
rlabel metal4 s 25270 22104 25330 22304 4 ui_in[1]
port 7 nsew
rlabel metal4 s 24718 22104 24778 22304 4 ui_in[2]
port 8 nsew
rlabel metal4 s 24166 22104 24226 22304 4 ui_in[3]
port 9 nsew
rlabel metal4 s 23614 22104 23674 22304 4 ui_in[4]
port 10 nsew
rlabel metal4 s 23062 22104 23122 22304 4 ui_in[5]
port 11 nsew
rlabel metal4 s 22510 22104 22570 22304 4 ui_in[6]
port 12 nsew
rlabel metal4 s 21958 22104 22018 22304 4 ui_in[7]
port 13 nsew
rlabel metal4 s 21406 22104 21466 22304 4 uio_in[0]
port 14 nsew
rlabel metal4 s 20854 22104 20914 22304 4 uio_in[1]
port 15 nsew
rlabel metal4 s 20302 22104 20362 22304 4 uio_in[2]
port 16 nsew
rlabel metal4 s 19750 22104 19810 22304 4 uio_in[3]
port 17 nsew
rlabel metal4 s 19198 22104 19258 22304 4 uio_in[4]
port 18 nsew
rlabel metal4 s 18646 22104 18706 22304 4 uio_in[5]
port 19 nsew
rlabel metal4 s 18094 22104 18154 22304 4 uio_in[6]
port 20 nsew
rlabel metal4 s 17542 22104 17602 22304 4 uio_in[7]
port 21 nsew
rlabel metal4 s 8158 22104 8218 22304 4 uio_oe[0]
port 22 nsew
rlabel metal4 s 7606 22104 7666 22304 4 uio_oe[1]
port 23 nsew
rlabel metal4 s 7054 22104 7114 22304 4 uio_oe[2]
port 24 nsew
rlabel metal4 s 6502 22104 6562 22304 4 uio_oe[3]
port 25 nsew
rlabel metal4 s 5950 22104 6010 22304 4 uio_oe[4]
port 26 nsew
rlabel metal4 s 5398 22104 5458 22304 4 uio_oe[5]
port 27 nsew
rlabel metal4 s 4846 22104 4906 22304 4 uio_oe[6]
port 28 nsew
rlabel metal4 s 4294 22104 4354 22304 4 uio_oe[7]
port 29 nsew
rlabel metal4 s 12574 22104 12634 22304 4 uio_out[0]
port 30 nsew
rlabel metal4 s 12022 22104 12082 22304 4 uio_out[1]
port 31 nsew
rlabel metal4 s 11470 22104 11530 22304 4 uio_out[2]
port 32 nsew
rlabel metal4 s 10918 22104 10978 22304 4 uio_out[3]
port 33 nsew
rlabel metal4 s 10366 22104 10426 22304 4 uio_out[4]
port 34 nsew
rlabel metal4 s 9814 22104 9874 22304 4 uio_out[5]
port 35 nsew
rlabel metal4 s 9262 22104 9322 22304 4 uio_out[6]
port 36 nsew
rlabel metal4 s 8710 22104 8770 22304 4 uio_out[7]
port 37 nsew
rlabel metal4 s 16990 22104 17050 22304 4 uo_out[0]
port 38 nsew
rlabel metal4 s 16438 22104 16498 22304 4 uo_out[1]
port 39 nsew
rlabel metal4 s 15886 22104 15946 22304 4 uo_out[2]
port 40 nsew
rlabel metal4 s 15334 22104 15394 22304 4 uo_out[3]
port 41 nsew
rlabel metal4 s 14782 22104 14842 22304 4 uo_out[4]
port 42 nsew
rlabel metal4 s 14230 22104 14290 22304 4 uo_out[5]
port 43 nsew
rlabel metal4 s 13678 22104 13738 22304 4 uo_out[6]
port 44 nsew
rlabel metal4 s 13126 22104 13186 22304 4 uo_out[7]
port 45 nsew
flabel metal4 s 0 0 400 22304 0 FreeSans 2000 0 0 0 VPWR
port 46 nsew
<< end >>
