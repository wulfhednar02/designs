magic
tech sky130A
magscale 1 2
timestamp 1699066547
<< error_s >>
rect 3385 516 3397 522
rect 3407 516 3419 522
rect 3373 498 3375 510
rect 3430 498 3431 510
rect 116 372 122 378
rect 146 348 152 368
rect 188 260 194 280
rect 146 238 152 244
rect 3373 130 3375 142
rect 3430 130 3431 142
rect 3385 118 3397 124
rect 3407 118 3419 124
<< locali >>
rect 0 300 64 319
rect 0 266 7 300
rect 41 266 64 300
rect 0 245 64 266
rect 302 263 347 303
rect 1228 263 1440 303
<< viali >>
rect 3385 476 3419 510
rect 3385 390 3419 424
rect 3385 303 3419 337
rect 7 266 41 300
rect 86 266 120 300
rect 3385 216 3419 250
rect 3385 130 3419 164
<< metal1 >>
rect 3375 510 3430 516
rect 3375 476 3385 510
rect 3419 476 3430 510
rect 3375 424 3430 476
rect 3375 390 3385 424
rect 3419 390 3430 424
rect 3375 337 3430 390
rect 0 300 132 319
rect 0 266 7 300
rect 41 266 86 300
rect 120 266 132 300
rect 0 245 132 266
rect 3375 303 3385 337
rect 3419 303 3430 337
rect 3375 250 3430 303
rect 3375 216 3385 250
rect 3419 216 3430 250
rect 3375 164 3430 216
rect 3375 130 3385 164
rect 3419 130 3430 164
rect 3375 124 3430 130
<< via1 >>
rect 63 566 115 618
rect 155 566 207 618
rect 247 566 299 618
rect 339 566 391 618
rect 431 566 483 618
rect 523 566 575 618
rect 615 566 667 618
rect 707 566 759 618
rect 799 566 851 618
rect 891 566 943 618
rect 983 566 1035 618
rect 1075 566 1127 618
rect 1167 566 1219 618
rect 1259 566 1311 618
rect 1351 566 1403 618
rect 1443 566 1495 618
rect 1535 566 1587 618
rect 1627 566 1679 618
rect 1719 566 1771 618
rect 1811 566 1863 618
rect 1903 566 1955 618
rect 1995 566 2047 618
rect 2087 566 2139 618
rect 2179 566 2231 618
rect 2271 566 2323 618
rect 2363 566 2415 618
rect 2455 566 2507 618
rect 2547 566 2599 618
rect 2639 566 2691 618
rect 2731 566 2783 618
rect 2823 566 2875 618
rect 2915 566 2967 618
rect 3007 566 3059 618
rect 3099 566 3151 618
rect 3191 566 3243 618
rect 3283 566 3335 618
rect 3375 566 3427 618
rect 63 22 115 74
rect 155 22 207 74
rect 247 22 299 74
rect 339 22 391 74
rect 431 22 483 74
rect 523 22 575 74
rect 615 22 667 74
rect 707 22 759 74
rect 799 22 851 74
rect 891 22 943 74
rect 983 22 1035 74
rect 1075 22 1127 74
rect 1167 22 1219 74
rect 1259 22 1311 74
rect 1351 22 1403 74
rect 1443 22 1495 74
rect 1535 22 1587 74
rect 1627 22 1679 74
rect 1719 22 1771 74
rect 1811 22 1863 74
rect 1903 22 1955 74
rect 1995 22 2047 74
rect 2087 22 2139 74
rect 2179 22 2231 74
rect 2271 22 2323 74
rect 2363 22 2415 74
rect 2455 22 2507 74
rect 2547 22 2599 74
rect 2639 22 2691 74
rect 2731 22 2783 74
rect 2823 22 2875 74
rect 2915 22 2967 74
rect 3007 22 3059 74
rect 3099 22 3151 74
rect 3191 22 3243 74
rect 3283 22 3335 74
rect 3375 22 3427 74
<< metal2 >>
rect 43 618 3447 640
rect 43 566 63 618
rect 115 566 155 618
rect 207 566 247 618
rect 299 566 339 618
rect 391 566 431 618
rect 483 566 523 618
rect 575 566 615 618
rect 667 566 707 618
rect 759 566 799 618
rect 851 566 891 618
rect 943 566 983 618
rect 1035 566 1075 618
rect 1127 566 1167 618
rect 1219 566 1259 618
rect 1311 566 1351 618
rect 1403 566 1443 618
rect 1495 566 1535 618
rect 1587 566 1627 618
rect 1679 566 1719 618
rect 1771 566 1811 618
rect 1863 566 1903 618
rect 1955 566 1995 618
rect 2047 566 2087 618
rect 2139 566 2179 618
rect 2231 566 2271 618
rect 2323 566 2363 618
rect 2415 566 2455 618
rect 2507 566 2547 618
rect 2599 566 2639 618
rect 2691 566 2731 618
rect 2783 566 2823 618
rect 2875 566 2915 618
rect 2967 566 3007 618
rect 3059 566 3099 618
rect 3151 566 3191 618
rect 3243 566 3283 618
rect 3335 566 3375 618
rect 3427 566 3447 618
rect 43 544 3447 566
rect 43 74 3447 96
rect 43 22 63 74
rect 115 22 155 74
rect 207 22 247 74
rect 299 22 339 74
rect 391 22 431 74
rect 483 22 523 74
rect 575 22 615 74
rect 667 22 707 74
rect 759 22 799 74
rect 851 22 891 74
rect 943 22 983 74
rect 1035 22 1075 74
rect 1127 22 1167 74
rect 1219 22 1259 74
rect 1311 22 1351 74
rect 1403 22 1443 74
rect 1495 22 1535 74
rect 1587 22 1627 74
rect 1679 22 1719 74
rect 1771 22 1811 74
rect 1863 22 1903 74
rect 1955 22 1995 74
rect 2047 22 2087 74
rect 2139 22 2179 74
rect 2231 22 2271 74
rect 2323 22 2363 74
rect 2415 22 2455 74
rect 2507 22 2547 74
rect 2599 22 2639 74
rect 2691 22 2731 74
rect 2783 22 2823 74
rect 2875 22 2915 74
rect 2967 22 3007 74
rect 3059 22 3099 74
rect 3151 22 3191 74
rect 3243 22 3283 74
rect 3335 22 3375 74
rect 3427 22 3447 74
rect 43 0 3447 22
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1699066547
transform 1 0 43 0 1 48
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_0
timestamp 1699066547
transform 1 0 319 0 1 48
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_0
timestamp 1699066547
transform 1 0 1423 0 1 48
box -38 -48 2062 592
<< labels >>
flabel metal1 s 0 245 132 319 0 FreeSans 224 0 0 0 IN
port 2 nsew
flabel metal1 s 3375 126 3430 515 0 FreeSans 44 0 0 0 OUT
port 3 nsew
flabel metal1 s 3402 142 3402 142 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 3403 320 3403 320 0 FreeSans 44 0 0 0 OUT
flabel metal2 s 43 0 3447 96 0 FreeSans 44 0 0 0 VSS
port 5 nsew
flabel metal2 s 3408 50 3408 50 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 1734 53 1734 53 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 787 50 787 50 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 2655 57 2655 57 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 43 544 3447 640 0 FreeSans 44 0 0 0 VDD
port 6 nsew
flabel metal2 s 3395 598 3395 598 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 1732 596 1732 596 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 796 594 796 594 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 2675 596 2675 596 0 FreeSans 44 0 0 0 VDD
<< end >>
