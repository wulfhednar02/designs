magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< nwell >>
rect -61 -76 1534 8144
<< pmos >>
rect 204 0 1004 8000
<< pdiff >>
rect 0 7977 204 8000
rect 0 7943 13 7977
rect 47 7943 85 7977
rect 119 7943 157 7977
rect 191 7943 204 7977
rect 0 7905 204 7943
rect 0 7871 13 7905
rect 47 7871 85 7905
rect 119 7871 157 7905
rect 191 7871 204 7905
rect 0 7833 204 7871
rect 0 7799 13 7833
rect 47 7799 85 7833
rect 119 7799 157 7833
rect 191 7799 204 7833
rect 0 7761 204 7799
rect 0 7727 13 7761
rect 47 7727 85 7761
rect 119 7727 157 7761
rect 191 7727 204 7761
rect 0 7689 204 7727
rect 0 7655 13 7689
rect 47 7655 85 7689
rect 119 7655 157 7689
rect 191 7655 204 7689
rect 0 7617 204 7655
rect 0 7583 13 7617
rect 47 7583 85 7617
rect 119 7583 157 7617
rect 191 7583 204 7617
rect 0 7545 204 7583
rect 0 7511 13 7545
rect 47 7511 85 7545
rect 119 7511 157 7545
rect 191 7511 204 7545
rect 0 7473 204 7511
rect 0 7439 13 7473
rect 47 7439 85 7473
rect 119 7439 157 7473
rect 191 7439 204 7473
rect 0 7401 204 7439
rect 0 7367 13 7401
rect 47 7367 85 7401
rect 119 7367 157 7401
rect 191 7367 204 7401
rect 0 7329 204 7367
rect 0 7295 13 7329
rect 47 7295 85 7329
rect 119 7295 157 7329
rect 191 7295 204 7329
rect 0 7257 204 7295
rect 0 7223 13 7257
rect 47 7223 85 7257
rect 119 7223 157 7257
rect 191 7223 204 7257
rect 0 7185 204 7223
rect 0 7151 13 7185
rect 47 7151 85 7185
rect 119 7151 157 7185
rect 191 7151 204 7185
rect 0 7113 204 7151
rect 0 7079 13 7113
rect 47 7079 85 7113
rect 119 7079 157 7113
rect 191 7079 204 7113
rect 0 7041 204 7079
rect 0 7007 13 7041
rect 47 7007 85 7041
rect 119 7007 157 7041
rect 191 7007 204 7041
rect 0 6969 204 7007
rect 0 6935 13 6969
rect 47 6935 85 6969
rect 119 6935 157 6969
rect 191 6935 204 6969
rect 0 6897 204 6935
rect 0 6863 13 6897
rect 47 6863 85 6897
rect 119 6863 157 6897
rect 191 6863 204 6897
rect 0 6825 204 6863
rect 0 6791 13 6825
rect 47 6791 85 6825
rect 119 6791 157 6825
rect 191 6791 204 6825
rect 0 6753 204 6791
rect 0 6719 13 6753
rect 47 6719 85 6753
rect 119 6719 157 6753
rect 191 6719 204 6753
rect 0 6681 204 6719
rect 0 6647 13 6681
rect 47 6647 85 6681
rect 119 6647 157 6681
rect 191 6647 204 6681
rect 0 6609 204 6647
rect 0 6575 13 6609
rect 47 6575 85 6609
rect 119 6575 157 6609
rect 191 6575 204 6609
rect 0 6537 204 6575
rect 0 6503 13 6537
rect 47 6503 85 6537
rect 119 6503 157 6537
rect 191 6503 204 6537
rect 0 6465 204 6503
rect 0 6431 13 6465
rect 47 6431 85 6465
rect 119 6431 157 6465
rect 191 6431 204 6465
rect 0 6393 204 6431
rect 0 6359 13 6393
rect 47 6359 85 6393
rect 119 6359 157 6393
rect 191 6359 204 6393
rect 0 6321 204 6359
rect 0 6287 13 6321
rect 47 6287 85 6321
rect 119 6287 157 6321
rect 191 6287 204 6321
rect 0 6249 204 6287
rect 0 6215 13 6249
rect 47 6215 85 6249
rect 119 6215 157 6249
rect 191 6215 204 6249
rect 0 6177 204 6215
rect 0 6143 13 6177
rect 47 6143 85 6177
rect 119 6143 157 6177
rect 191 6143 204 6177
rect 0 6105 204 6143
rect 0 6071 13 6105
rect 47 6071 85 6105
rect 119 6071 157 6105
rect 191 6071 204 6105
rect 0 6033 204 6071
rect 0 5999 13 6033
rect 47 5999 85 6033
rect 119 5999 157 6033
rect 191 5999 204 6033
rect 0 5961 204 5999
rect 0 5927 13 5961
rect 47 5927 85 5961
rect 119 5927 157 5961
rect 191 5927 204 5961
rect 0 5889 204 5927
rect 0 5855 13 5889
rect 47 5855 85 5889
rect 119 5855 157 5889
rect 191 5855 204 5889
rect 0 5817 204 5855
rect 0 5783 13 5817
rect 47 5783 85 5817
rect 119 5783 157 5817
rect 191 5783 204 5817
rect 0 5745 204 5783
rect 0 5711 13 5745
rect 47 5711 85 5745
rect 119 5711 157 5745
rect 191 5711 204 5745
rect 0 5673 204 5711
rect 0 5639 13 5673
rect 47 5639 85 5673
rect 119 5639 157 5673
rect 191 5639 204 5673
rect 0 5601 204 5639
rect 0 5567 13 5601
rect 47 5567 85 5601
rect 119 5567 157 5601
rect 191 5567 204 5601
rect 0 5529 204 5567
rect 0 5495 13 5529
rect 47 5495 85 5529
rect 119 5495 157 5529
rect 191 5495 204 5529
rect 0 5457 204 5495
rect 0 5423 13 5457
rect 47 5423 85 5457
rect 119 5423 157 5457
rect 191 5423 204 5457
rect 0 5385 204 5423
rect 0 5351 13 5385
rect 47 5351 85 5385
rect 119 5351 157 5385
rect 191 5351 204 5385
rect 0 5313 204 5351
rect 0 5279 13 5313
rect 47 5279 85 5313
rect 119 5279 157 5313
rect 191 5279 204 5313
rect 0 5241 204 5279
rect 0 5207 13 5241
rect 47 5207 85 5241
rect 119 5207 157 5241
rect 191 5207 204 5241
rect 0 5169 204 5207
rect 0 5135 13 5169
rect 47 5135 85 5169
rect 119 5135 157 5169
rect 191 5135 204 5169
rect 0 5097 204 5135
rect 0 5063 13 5097
rect 47 5063 85 5097
rect 119 5063 157 5097
rect 191 5063 204 5097
rect 0 5025 204 5063
rect 0 4991 13 5025
rect 47 4991 85 5025
rect 119 4991 157 5025
rect 191 4991 204 5025
rect 0 4953 204 4991
rect 0 4919 13 4953
rect 47 4919 85 4953
rect 119 4919 157 4953
rect 191 4919 204 4953
rect 0 4881 204 4919
rect 0 4847 13 4881
rect 47 4847 85 4881
rect 119 4847 157 4881
rect 191 4847 204 4881
rect 0 4809 204 4847
rect 0 4775 13 4809
rect 47 4775 85 4809
rect 119 4775 157 4809
rect 191 4775 204 4809
rect 0 4737 204 4775
rect 0 4703 13 4737
rect 47 4703 85 4737
rect 119 4703 157 4737
rect 191 4703 204 4737
rect 0 4665 204 4703
rect 0 4631 13 4665
rect 47 4631 85 4665
rect 119 4631 157 4665
rect 191 4631 204 4665
rect 0 4593 204 4631
rect 0 4559 13 4593
rect 47 4559 85 4593
rect 119 4559 157 4593
rect 191 4559 204 4593
rect 0 4521 204 4559
rect 0 4487 13 4521
rect 47 4487 85 4521
rect 119 4487 157 4521
rect 191 4487 204 4521
rect 0 4449 204 4487
rect 0 4415 13 4449
rect 47 4415 85 4449
rect 119 4415 157 4449
rect 191 4415 204 4449
rect 0 4377 204 4415
rect 0 4343 13 4377
rect 47 4343 85 4377
rect 119 4343 157 4377
rect 191 4343 204 4377
rect 0 4305 204 4343
rect 0 4271 13 4305
rect 47 4271 85 4305
rect 119 4271 157 4305
rect 191 4271 204 4305
rect 0 4233 204 4271
rect 0 4199 13 4233
rect 47 4199 85 4233
rect 119 4199 157 4233
rect 191 4199 204 4233
rect 0 4161 204 4199
rect 0 4127 13 4161
rect 47 4127 85 4161
rect 119 4127 157 4161
rect 191 4127 204 4161
rect 0 4089 204 4127
rect 0 4055 13 4089
rect 47 4055 85 4089
rect 119 4055 157 4089
rect 191 4055 204 4089
rect 0 4017 204 4055
rect 0 3983 13 4017
rect 47 3983 85 4017
rect 119 3983 157 4017
rect 191 3983 204 4017
rect 0 3945 204 3983
rect 0 3911 13 3945
rect 47 3911 85 3945
rect 119 3911 157 3945
rect 191 3911 204 3945
rect 0 3873 204 3911
rect 0 3839 13 3873
rect 47 3839 85 3873
rect 119 3839 157 3873
rect 191 3839 204 3873
rect 0 3801 204 3839
rect 0 3767 13 3801
rect 47 3767 85 3801
rect 119 3767 157 3801
rect 191 3767 204 3801
rect 0 3729 204 3767
rect 0 3695 13 3729
rect 47 3695 85 3729
rect 119 3695 157 3729
rect 191 3695 204 3729
rect 0 3657 204 3695
rect 0 3623 13 3657
rect 47 3623 85 3657
rect 119 3623 157 3657
rect 191 3623 204 3657
rect 0 3585 204 3623
rect 0 3551 13 3585
rect 47 3551 85 3585
rect 119 3551 157 3585
rect 191 3551 204 3585
rect 0 3513 204 3551
rect 0 3479 13 3513
rect 47 3479 85 3513
rect 119 3479 157 3513
rect 191 3479 204 3513
rect 0 3441 204 3479
rect 0 3407 13 3441
rect 47 3407 85 3441
rect 119 3407 157 3441
rect 191 3407 204 3441
rect 0 3369 204 3407
rect 0 3335 13 3369
rect 47 3335 85 3369
rect 119 3335 157 3369
rect 191 3335 204 3369
rect 0 3297 204 3335
rect 0 3263 13 3297
rect 47 3263 85 3297
rect 119 3263 157 3297
rect 191 3263 204 3297
rect 0 3225 204 3263
rect 0 3191 13 3225
rect 47 3191 85 3225
rect 119 3191 157 3225
rect 191 3191 204 3225
rect 0 3153 204 3191
rect 0 3119 13 3153
rect 47 3119 85 3153
rect 119 3119 157 3153
rect 191 3119 204 3153
rect 0 3081 204 3119
rect 0 3047 13 3081
rect 47 3047 85 3081
rect 119 3047 157 3081
rect 191 3047 204 3081
rect 0 3009 204 3047
rect 0 2975 13 3009
rect 47 2975 85 3009
rect 119 2975 157 3009
rect 191 2975 204 3009
rect 0 2937 204 2975
rect 0 2903 13 2937
rect 47 2903 85 2937
rect 119 2903 157 2937
rect 191 2903 204 2937
rect 0 2865 204 2903
rect 0 2831 13 2865
rect 47 2831 85 2865
rect 119 2831 157 2865
rect 191 2831 204 2865
rect 0 2793 204 2831
rect 0 2759 13 2793
rect 47 2759 85 2793
rect 119 2759 157 2793
rect 191 2759 204 2793
rect 0 2721 204 2759
rect 0 2687 13 2721
rect 47 2687 85 2721
rect 119 2687 157 2721
rect 191 2687 204 2721
rect 0 2649 204 2687
rect 0 2615 13 2649
rect 47 2615 85 2649
rect 119 2615 157 2649
rect 191 2615 204 2649
rect 0 2577 204 2615
rect 0 2543 13 2577
rect 47 2543 85 2577
rect 119 2543 157 2577
rect 191 2543 204 2577
rect 0 2505 204 2543
rect 0 2471 13 2505
rect 47 2471 85 2505
rect 119 2471 157 2505
rect 191 2471 204 2505
rect 0 2433 204 2471
rect 0 2399 13 2433
rect 47 2399 85 2433
rect 119 2399 157 2433
rect 191 2399 204 2433
rect 0 2361 204 2399
rect 0 2327 13 2361
rect 47 2327 85 2361
rect 119 2327 157 2361
rect 191 2327 204 2361
rect 0 2289 204 2327
rect 0 2255 13 2289
rect 47 2255 85 2289
rect 119 2255 157 2289
rect 191 2255 204 2289
rect 0 2217 204 2255
rect 0 2183 13 2217
rect 47 2183 85 2217
rect 119 2183 157 2217
rect 191 2183 204 2217
rect 0 2145 204 2183
rect 0 2111 13 2145
rect 47 2111 85 2145
rect 119 2111 157 2145
rect 191 2111 204 2145
rect 0 2073 204 2111
rect 0 2039 13 2073
rect 47 2039 85 2073
rect 119 2039 157 2073
rect 191 2039 204 2073
rect 0 2001 204 2039
rect 0 1967 13 2001
rect 47 1967 85 2001
rect 119 1967 157 2001
rect 191 1967 204 2001
rect 0 1929 204 1967
rect 0 1895 13 1929
rect 47 1895 85 1929
rect 119 1895 157 1929
rect 191 1895 204 1929
rect 0 1857 204 1895
rect 0 1823 13 1857
rect 47 1823 85 1857
rect 119 1823 157 1857
rect 191 1823 204 1857
rect 0 1785 204 1823
rect 0 1751 13 1785
rect 47 1751 85 1785
rect 119 1751 157 1785
rect 191 1751 204 1785
rect 0 1713 204 1751
rect 0 1679 13 1713
rect 47 1679 85 1713
rect 119 1679 157 1713
rect 191 1679 204 1713
rect 0 1641 204 1679
rect 0 1607 13 1641
rect 47 1607 85 1641
rect 119 1607 157 1641
rect 191 1607 204 1641
rect 0 1569 204 1607
rect 0 1535 13 1569
rect 47 1535 85 1569
rect 119 1535 157 1569
rect 191 1535 204 1569
rect 0 1497 204 1535
rect 0 1463 13 1497
rect 47 1463 85 1497
rect 119 1463 157 1497
rect 191 1463 204 1497
rect 0 1425 204 1463
rect 0 1391 13 1425
rect 47 1391 85 1425
rect 119 1391 157 1425
rect 191 1391 204 1425
rect 0 1353 204 1391
rect 0 1319 13 1353
rect 47 1319 85 1353
rect 119 1319 157 1353
rect 191 1319 204 1353
rect 0 1281 204 1319
rect 0 1247 13 1281
rect 47 1247 85 1281
rect 119 1247 157 1281
rect 191 1247 204 1281
rect 0 1209 204 1247
rect 0 1175 13 1209
rect 47 1175 85 1209
rect 119 1175 157 1209
rect 191 1175 204 1209
rect 0 1137 204 1175
rect 0 1103 13 1137
rect 47 1103 85 1137
rect 119 1103 157 1137
rect 191 1103 204 1137
rect 0 1065 204 1103
rect 0 1031 13 1065
rect 47 1031 85 1065
rect 119 1031 157 1065
rect 191 1031 204 1065
rect 0 993 204 1031
rect 0 959 13 993
rect 47 959 85 993
rect 119 959 157 993
rect 191 959 204 993
rect 0 921 204 959
rect 0 887 13 921
rect 47 887 85 921
rect 119 887 157 921
rect 191 887 204 921
rect 0 849 204 887
rect 0 815 13 849
rect 47 815 85 849
rect 119 815 157 849
rect 191 815 204 849
rect 0 777 204 815
rect 0 743 13 777
rect 47 743 85 777
rect 119 743 157 777
rect 191 743 204 777
rect 0 705 204 743
rect 0 671 13 705
rect 47 671 85 705
rect 119 671 157 705
rect 191 671 204 705
rect 0 633 204 671
rect 0 599 13 633
rect 47 599 85 633
rect 119 599 157 633
rect 191 599 204 633
rect 0 561 204 599
rect 0 527 13 561
rect 47 527 85 561
rect 119 527 157 561
rect 191 527 204 561
rect 0 489 204 527
rect 0 455 13 489
rect 47 455 85 489
rect 119 455 157 489
rect 191 455 204 489
rect 0 417 204 455
rect 0 383 13 417
rect 47 383 85 417
rect 119 383 157 417
rect 191 383 204 417
rect 0 345 204 383
rect 0 311 13 345
rect 47 311 85 345
rect 119 311 157 345
rect 191 311 204 345
rect 0 273 204 311
rect 0 239 13 273
rect 47 239 85 273
rect 119 239 157 273
rect 191 239 204 273
rect 0 201 204 239
rect 0 167 13 201
rect 47 167 85 201
rect 119 167 157 201
rect 191 167 204 201
rect 0 129 204 167
rect 0 95 13 129
rect 47 95 85 129
rect 119 95 157 129
rect 191 95 204 129
rect 0 57 204 95
rect 0 23 13 57
rect 47 23 85 57
rect 119 23 157 57
rect 191 23 204 57
rect 0 0 204 23
rect 1004 7977 1208 8000
rect 1004 7943 1017 7977
rect 1051 7943 1089 7977
rect 1123 7943 1161 7977
rect 1195 7943 1208 7977
rect 1004 7905 1208 7943
rect 1004 7871 1017 7905
rect 1051 7871 1089 7905
rect 1123 7871 1161 7905
rect 1195 7871 1208 7905
rect 1004 7833 1208 7871
rect 1004 7799 1017 7833
rect 1051 7799 1089 7833
rect 1123 7799 1161 7833
rect 1195 7799 1208 7833
rect 1004 7761 1208 7799
rect 1004 7727 1017 7761
rect 1051 7727 1089 7761
rect 1123 7727 1161 7761
rect 1195 7727 1208 7761
rect 1004 7689 1208 7727
rect 1004 7655 1017 7689
rect 1051 7655 1089 7689
rect 1123 7655 1161 7689
rect 1195 7655 1208 7689
rect 1004 7617 1208 7655
rect 1004 7583 1017 7617
rect 1051 7583 1089 7617
rect 1123 7583 1161 7617
rect 1195 7583 1208 7617
rect 1004 7545 1208 7583
rect 1004 7511 1017 7545
rect 1051 7511 1089 7545
rect 1123 7511 1161 7545
rect 1195 7511 1208 7545
rect 1004 7473 1208 7511
rect 1004 7439 1017 7473
rect 1051 7439 1089 7473
rect 1123 7439 1161 7473
rect 1195 7439 1208 7473
rect 1004 7401 1208 7439
rect 1004 7367 1017 7401
rect 1051 7367 1089 7401
rect 1123 7367 1161 7401
rect 1195 7367 1208 7401
rect 1004 7329 1208 7367
rect 1004 7295 1017 7329
rect 1051 7295 1089 7329
rect 1123 7295 1161 7329
rect 1195 7295 1208 7329
rect 1004 7257 1208 7295
rect 1004 7223 1017 7257
rect 1051 7223 1089 7257
rect 1123 7223 1161 7257
rect 1195 7223 1208 7257
rect 1004 7185 1208 7223
rect 1004 7151 1017 7185
rect 1051 7151 1089 7185
rect 1123 7151 1161 7185
rect 1195 7151 1208 7185
rect 1004 7113 1208 7151
rect 1004 7079 1017 7113
rect 1051 7079 1089 7113
rect 1123 7079 1161 7113
rect 1195 7079 1208 7113
rect 1004 7041 1208 7079
rect 1004 7007 1017 7041
rect 1051 7007 1089 7041
rect 1123 7007 1161 7041
rect 1195 7007 1208 7041
rect 1004 6969 1208 7007
rect 1004 6935 1017 6969
rect 1051 6935 1089 6969
rect 1123 6935 1161 6969
rect 1195 6935 1208 6969
rect 1004 6897 1208 6935
rect 1004 6863 1017 6897
rect 1051 6863 1089 6897
rect 1123 6863 1161 6897
rect 1195 6863 1208 6897
rect 1004 6825 1208 6863
rect 1004 6791 1017 6825
rect 1051 6791 1089 6825
rect 1123 6791 1161 6825
rect 1195 6791 1208 6825
rect 1004 6753 1208 6791
rect 1004 6719 1017 6753
rect 1051 6719 1089 6753
rect 1123 6719 1161 6753
rect 1195 6719 1208 6753
rect 1004 6681 1208 6719
rect 1004 6647 1017 6681
rect 1051 6647 1089 6681
rect 1123 6647 1161 6681
rect 1195 6647 1208 6681
rect 1004 6609 1208 6647
rect 1004 6575 1017 6609
rect 1051 6575 1089 6609
rect 1123 6575 1161 6609
rect 1195 6575 1208 6609
rect 1004 6537 1208 6575
rect 1004 6503 1017 6537
rect 1051 6503 1089 6537
rect 1123 6503 1161 6537
rect 1195 6503 1208 6537
rect 1004 6465 1208 6503
rect 1004 6431 1017 6465
rect 1051 6431 1089 6465
rect 1123 6431 1161 6465
rect 1195 6431 1208 6465
rect 1004 6393 1208 6431
rect 1004 6359 1017 6393
rect 1051 6359 1089 6393
rect 1123 6359 1161 6393
rect 1195 6359 1208 6393
rect 1004 6321 1208 6359
rect 1004 6287 1017 6321
rect 1051 6287 1089 6321
rect 1123 6287 1161 6321
rect 1195 6287 1208 6321
rect 1004 6249 1208 6287
rect 1004 6215 1017 6249
rect 1051 6215 1089 6249
rect 1123 6215 1161 6249
rect 1195 6215 1208 6249
rect 1004 6177 1208 6215
rect 1004 6143 1017 6177
rect 1051 6143 1089 6177
rect 1123 6143 1161 6177
rect 1195 6143 1208 6177
rect 1004 6105 1208 6143
rect 1004 6071 1017 6105
rect 1051 6071 1089 6105
rect 1123 6071 1161 6105
rect 1195 6071 1208 6105
rect 1004 6033 1208 6071
rect 1004 5999 1017 6033
rect 1051 5999 1089 6033
rect 1123 5999 1161 6033
rect 1195 5999 1208 6033
rect 1004 5961 1208 5999
rect 1004 5927 1017 5961
rect 1051 5927 1089 5961
rect 1123 5927 1161 5961
rect 1195 5927 1208 5961
rect 1004 5889 1208 5927
rect 1004 5855 1017 5889
rect 1051 5855 1089 5889
rect 1123 5855 1161 5889
rect 1195 5855 1208 5889
rect 1004 5817 1208 5855
rect 1004 5783 1017 5817
rect 1051 5783 1089 5817
rect 1123 5783 1161 5817
rect 1195 5783 1208 5817
rect 1004 5745 1208 5783
rect 1004 5711 1017 5745
rect 1051 5711 1089 5745
rect 1123 5711 1161 5745
rect 1195 5711 1208 5745
rect 1004 5673 1208 5711
rect 1004 5639 1017 5673
rect 1051 5639 1089 5673
rect 1123 5639 1161 5673
rect 1195 5639 1208 5673
rect 1004 5601 1208 5639
rect 1004 5567 1017 5601
rect 1051 5567 1089 5601
rect 1123 5567 1161 5601
rect 1195 5567 1208 5601
rect 1004 5529 1208 5567
rect 1004 5495 1017 5529
rect 1051 5495 1089 5529
rect 1123 5495 1161 5529
rect 1195 5495 1208 5529
rect 1004 5457 1208 5495
rect 1004 5423 1017 5457
rect 1051 5423 1089 5457
rect 1123 5423 1161 5457
rect 1195 5423 1208 5457
rect 1004 5385 1208 5423
rect 1004 5351 1017 5385
rect 1051 5351 1089 5385
rect 1123 5351 1161 5385
rect 1195 5351 1208 5385
rect 1004 5313 1208 5351
rect 1004 5279 1017 5313
rect 1051 5279 1089 5313
rect 1123 5279 1161 5313
rect 1195 5279 1208 5313
rect 1004 5241 1208 5279
rect 1004 5207 1017 5241
rect 1051 5207 1089 5241
rect 1123 5207 1161 5241
rect 1195 5207 1208 5241
rect 1004 5169 1208 5207
rect 1004 5135 1017 5169
rect 1051 5135 1089 5169
rect 1123 5135 1161 5169
rect 1195 5135 1208 5169
rect 1004 5097 1208 5135
rect 1004 5063 1017 5097
rect 1051 5063 1089 5097
rect 1123 5063 1161 5097
rect 1195 5063 1208 5097
rect 1004 5025 1208 5063
rect 1004 4991 1017 5025
rect 1051 4991 1089 5025
rect 1123 4991 1161 5025
rect 1195 4991 1208 5025
rect 1004 4953 1208 4991
rect 1004 4919 1017 4953
rect 1051 4919 1089 4953
rect 1123 4919 1161 4953
rect 1195 4919 1208 4953
rect 1004 4881 1208 4919
rect 1004 4847 1017 4881
rect 1051 4847 1089 4881
rect 1123 4847 1161 4881
rect 1195 4847 1208 4881
rect 1004 4809 1208 4847
rect 1004 4775 1017 4809
rect 1051 4775 1089 4809
rect 1123 4775 1161 4809
rect 1195 4775 1208 4809
rect 1004 4737 1208 4775
rect 1004 4703 1017 4737
rect 1051 4703 1089 4737
rect 1123 4703 1161 4737
rect 1195 4703 1208 4737
rect 1004 4665 1208 4703
rect 1004 4631 1017 4665
rect 1051 4631 1089 4665
rect 1123 4631 1161 4665
rect 1195 4631 1208 4665
rect 1004 4593 1208 4631
rect 1004 4559 1017 4593
rect 1051 4559 1089 4593
rect 1123 4559 1161 4593
rect 1195 4559 1208 4593
rect 1004 4521 1208 4559
rect 1004 4487 1017 4521
rect 1051 4487 1089 4521
rect 1123 4487 1161 4521
rect 1195 4487 1208 4521
rect 1004 4449 1208 4487
rect 1004 4415 1017 4449
rect 1051 4415 1089 4449
rect 1123 4415 1161 4449
rect 1195 4415 1208 4449
rect 1004 4377 1208 4415
rect 1004 4343 1017 4377
rect 1051 4343 1089 4377
rect 1123 4343 1161 4377
rect 1195 4343 1208 4377
rect 1004 4305 1208 4343
rect 1004 4271 1017 4305
rect 1051 4271 1089 4305
rect 1123 4271 1161 4305
rect 1195 4271 1208 4305
rect 1004 4233 1208 4271
rect 1004 4199 1017 4233
rect 1051 4199 1089 4233
rect 1123 4199 1161 4233
rect 1195 4199 1208 4233
rect 1004 4161 1208 4199
rect 1004 4127 1017 4161
rect 1051 4127 1089 4161
rect 1123 4127 1161 4161
rect 1195 4127 1208 4161
rect 1004 4089 1208 4127
rect 1004 4055 1017 4089
rect 1051 4055 1089 4089
rect 1123 4055 1161 4089
rect 1195 4055 1208 4089
rect 1004 4017 1208 4055
rect 1004 3983 1017 4017
rect 1051 3983 1089 4017
rect 1123 3983 1161 4017
rect 1195 3983 1208 4017
rect 1004 3945 1208 3983
rect 1004 3911 1017 3945
rect 1051 3911 1089 3945
rect 1123 3911 1161 3945
rect 1195 3911 1208 3945
rect 1004 3873 1208 3911
rect 1004 3839 1017 3873
rect 1051 3839 1089 3873
rect 1123 3839 1161 3873
rect 1195 3839 1208 3873
rect 1004 3801 1208 3839
rect 1004 3767 1017 3801
rect 1051 3767 1089 3801
rect 1123 3767 1161 3801
rect 1195 3767 1208 3801
rect 1004 3729 1208 3767
rect 1004 3695 1017 3729
rect 1051 3695 1089 3729
rect 1123 3695 1161 3729
rect 1195 3695 1208 3729
rect 1004 3657 1208 3695
rect 1004 3623 1017 3657
rect 1051 3623 1089 3657
rect 1123 3623 1161 3657
rect 1195 3623 1208 3657
rect 1004 3585 1208 3623
rect 1004 3551 1017 3585
rect 1051 3551 1089 3585
rect 1123 3551 1161 3585
rect 1195 3551 1208 3585
rect 1004 3513 1208 3551
rect 1004 3479 1017 3513
rect 1051 3479 1089 3513
rect 1123 3479 1161 3513
rect 1195 3479 1208 3513
rect 1004 3441 1208 3479
rect 1004 3407 1017 3441
rect 1051 3407 1089 3441
rect 1123 3407 1161 3441
rect 1195 3407 1208 3441
rect 1004 3369 1208 3407
rect 1004 3335 1017 3369
rect 1051 3335 1089 3369
rect 1123 3335 1161 3369
rect 1195 3335 1208 3369
rect 1004 3297 1208 3335
rect 1004 3263 1017 3297
rect 1051 3263 1089 3297
rect 1123 3263 1161 3297
rect 1195 3263 1208 3297
rect 1004 3225 1208 3263
rect 1004 3191 1017 3225
rect 1051 3191 1089 3225
rect 1123 3191 1161 3225
rect 1195 3191 1208 3225
rect 1004 3153 1208 3191
rect 1004 3119 1017 3153
rect 1051 3119 1089 3153
rect 1123 3119 1161 3153
rect 1195 3119 1208 3153
rect 1004 3081 1208 3119
rect 1004 3047 1017 3081
rect 1051 3047 1089 3081
rect 1123 3047 1161 3081
rect 1195 3047 1208 3081
rect 1004 3009 1208 3047
rect 1004 2975 1017 3009
rect 1051 2975 1089 3009
rect 1123 2975 1161 3009
rect 1195 2975 1208 3009
rect 1004 2937 1208 2975
rect 1004 2903 1017 2937
rect 1051 2903 1089 2937
rect 1123 2903 1161 2937
rect 1195 2903 1208 2937
rect 1004 2865 1208 2903
rect 1004 2831 1017 2865
rect 1051 2831 1089 2865
rect 1123 2831 1161 2865
rect 1195 2831 1208 2865
rect 1004 2793 1208 2831
rect 1004 2759 1017 2793
rect 1051 2759 1089 2793
rect 1123 2759 1161 2793
rect 1195 2759 1208 2793
rect 1004 2721 1208 2759
rect 1004 2687 1017 2721
rect 1051 2687 1089 2721
rect 1123 2687 1161 2721
rect 1195 2687 1208 2721
rect 1004 2649 1208 2687
rect 1004 2615 1017 2649
rect 1051 2615 1089 2649
rect 1123 2615 1161 2649
rect 1195 2615 1208 2649
rect 1004 2577 1208 2615
rect 1004 2543 1017 2577
rect 1051 2543 1089 2577
rect 1123 2543 1161 2577
rect 1195 2543 1208 2577
rect 1004 2505 1208 2543
rect 1004 2471 1017 2505
rect 1051 2471 1089 2505
rect 1123 2471 1161 2505
rect 1195 2471 1208 2505
rect 1004 2433 1208 2471
rect 1004 2399 1017 2433
rect 1051 2399 1089 2433
rect 1123 2399 1161 2433
rect 1195 2399 1208 2433
rect 1004 2361 1208 2399
rect 1004 2327 1017 2361
rect 1051 2327 1089 2361
rect 1123 2327 1161 2361
rect 1195 2327 1208 2361
rect 1004 2289 1208 2327
rect 1004 2255 1017 2289
rect 1051 2255 1089 2289
rect 1123 2255 1161 2289
rect 1195 2255 1208 2289
rect 1004 2217 1208 2255
rect 1004 2183 1017 2217
rect 1051 2183 1089 2217
rect 1123 2183 1161 2217
rect 1195 2183 1208 2217
rect 1004 2145 1208 2183
rect 1004 2111 1017 2145
rect 1051 2111 1089 2145
rect 1123 2111 1161 2145
rect 1195 2111 1208 2145
rect 1004 2073 1208 2111
rect 1004 2039 1017 2073
rect 1051 2039 1089 2073
rect 1123 2039 1161 2073
rect 1195 2039 1208 2073
rect 1004 2001 1208 2039
rect 1004 1967 1017 2001
rect 1051 1967 1089 2001
rect 1123 1967 1161 2001
rect 1195 1967 1208 2001
rect 1004 1929 1208 1967
rect 1004 1895 1017 1929
rect 1051 1895 1089 1929
rect 1123 1895 1161 1929
rect 1195 1895 1208 1929
rect 1004 1857 1208 1895
rect 1004 1823 1017 1857
rect 1051 1823 1089 1857
rect 1123 1823 1161 1857
rect 1195 1823 1208 1857
rect 1004 1785 1208 1823
rect 1004 1751 1017 1785
rect 1051 1751 1089 1785
rect 1123 1751 1161 1785
rect 1195 1751 1208 1785
rect 1004 1713 1208 1751
rect 1004 1679 1017 1713
rect 1051 1679 1089 1713
rect 1123 1679 1161 1713
rect 1195 1679 1208 1713
rect 1004 1641 1208 1679
rect 1004 1607 1017 1641
rect 1051 1607 1089 1641
rect 1123 1607 1161 1641
rect 1195 1607 1208 1641
rect 1004 1569 1208 1607
rect 1004 1535 1017 1569
rect 1051 1535 1089 1569
rect 1123 1535 1161 1569
rect 1195 1535 1208 1569
rect 1004 1497 1208 1535
rect 1004 1463 1017 1497
rect 1051 1463 1089 1497
rect 1123 1463 1161 1497
rect 1195 1463 1208 1497
rect 1004 1425 1208 1463
rect 1004 1391 1017 1425
rect 1051 1391 1089 1425
rect 1123 1391 1161 1425
rect 1195 1391 1208 1425
rect 1004 1353 1208 1391
rect 1004 1319 1017 1353
rect 1051 1319 1089 1353
rect 1123 1319 1161 1353
rect 1195 1319 1208 1353
rect 1004 1281 1208 1319
rect 1004 1247 1017 1281
rect 1051 1247 1089 1281
rect 1123 1247 1161 1281
rect 1195 1247 1208 1281
rect 1004 1209 1208 1247
rect 1004 1175 1017 1209
rect 1051 1175 1089 1209
rect 1123 1175 1161 1209
rect 1195 1175 1208 1209
rect 1004 1137 1208 1175
rect 1004 1103 1017 1137
rect 1051 1103 1089 1137
rect 1123 1103 1161 1137
rect 1195 1103 1208 1137
rect 1004 1065 1208 1103
rect 1004 1031 1017 1065
rect 1051 1031 1089 1065
rect 1123 1031 1161 1065
rect 1195 1031 1208 1065
rect 1004 993 1208 1031
rect 1004 959 1017 993
rect 1051 959 1089 993
rect 1123 959 1161 993
rect 1195 959 1208 993
rect 1004 921 1208 959
rect 1004 887 1017 921
rect 1051 887 1089 921
rect 1123 887 1161 921
rect 1195 887 1208 921
rect 1004 849 1208 887
rect 1004 815 1017 849
rect 1051 815 1089 849
rect 1123 815 1161 849
rect 1195 815 1208 849
rect 1004 777 1208 815
rect 1004 743 1017 777
rect 1051 743 1089 777
rect 1123 743 1161 777
rect 1195 743 1208 777
rect 1004 705 1208 743
rect 1004 671 1017 705
rect 1051 671 1089 705
rect 1123 671 1161 705
rect 1195 671 1208 705
rect 1004 633 1208 671
rect 1004 599 1017 633
rect 1051 599 1089 633
rect 1123 599 1161 633
rect 1195 599 1208 633
rect 1004 561 1208 599
rect 1004 527 1017 561
rect 1051 527 1089 561
rect 1123 527 1161 561
rect 1195 527 1208 561
rect 1004 489 1208 527
rect 1004 455 1017 489
rect 1051 455 1089 489
rect 1123 455 1161 489
rect 1195 455 1208 489
rect 1004 417 1208 455
rect 1004 383 1017 417
rect 1051 383 1089 417
rect 1123 383 1161 417
rect 1195 383 1208 417
rect 1004 345 1208 383
rect 1004 311 1017 345
rect 1051 311 1089 345
rect 1123 311 1161 345
rect 1195 311 1208 345
rect 1004 273 1208 311
rect 1004 239 1017 273
rect 1051 239 1089 273
rect 1123 239 1161 273
rect 1195 239 1208 273
rect 1004 201 1208 239
rect 1004 167 1017 201
rect 1051 167 1089 201
rect 1123 167 1161 201
rect 1195 167 1208 201
rect 1004 129 1208 167
rect 1004 95 1017 129
rect 1051 95 1089 129
rect 1123 95 1161 129
rect 1195 95 1208 129
rect 1004 57 1208 95
rect 1004 23 1017 57
rect 1051 23 1089 57
rect 1123 23 1161 57
rect 1195 23 1208 57
rect 1004 0 1208 23
<< pdiffc >>
rect 13 7943 47 7977
rect 85 7943 119 7977
rect 157 7943 191 7977
rect 13 7871 47 7905
rect 85 7871 119 7905
rect 157 7871 191 7905
rect 13 7799 47 7833
rect 85 7799 119 7833
rect 157 7799 191 7833
rect 13 7727 47 7761
rect 85 7727 119 7761
rect 157 7727 191 7761
rect 13 7655 47 7689
rect 85 7655 119 7689
rect 157 7655 191 7689
rect 13 7583 47 7617
rect 85 7583 119 7617
rect 157 7583 191 7617
rect 13 7511 47 7545
rect 85 7511 119 7545
rect 157 7511 191 7545
rect 13 7439 47 7473
rect 85 7439 119 7473
rect 157 7439 191 7473
rect 13 7367 47 7401
rect 85 7367 119 7401
rect 157 7367 191 7401
rect 13 7295 47 7329
rect 85 7295 119 7329
rect 157 7295 191 7329
rect 13 7223 47 7257
rect 85 7223 119 7257
rect 157 7223 191 7257
rect 13 7151 47 7185
rect 85 7151 119 7185
rect 157 7151 191 7185
rect 13 7079 47 7113
rect 85 7079 119 7113
rect 157 7079 191 7113
rect 13 7007 47 7041
rect 85 7007 119 7041
rect 157 7007 191 7041
rect 13 6935 47 6969
rect 85 6935 119 6969
rect 157 6935 191 6969
rect 13 6863 47 6897
rect 85 6863 119 6897
rect 157 6863 191 6897
rect 13 6791 47 6825
rect 85 6791 119 6825
rect 157 6791 191 6825
rect 13 6719 47 6753
rect 85 6719 119 6753
rect 157 6719 191 6753
rect 13 6647 47 6681
rect 85 6647 119 6681
rect 157 6647 191 6681
rect 13 6575 47 6609
rect 85 6575 119 6609
rect 157 6575 191 6609
rect 13 6503 47 6537
rect 85 6503 119 6537
rect 157 6503 191 6537
rect 13 6431 47 6465
rect 85 6431 119 6465
rect 157 6431 191 6465
rect 13 6359 47 6393
rect 85 6359 119 6393
rect 157 6359 191 6393
rect 13 6287 47 6321
rect 85 6287 119 6321
rect 157 6287 191 6321
rect 13 6215 47 6249
rect 85 6215 119 6249
rect 157 6215 191 6249
rect 13 6143 47 6177
rect 85 6143 119 6177
rect 157 6143 191 6177
rect 13 6071 47 6105
rect 85 6071 119 6105
rect 157 6071 191 6105
rect 13 5999 47 6033
rect 85 5999 119 6033
rect 157 5999 191 6033
rect 13 5927 47 5961
rect 85 5927 119 5961
rect 157 5927 191 5961
rect 13 5855 47 5889
rect 85 5855 119 5889
rect 157 5855 191 5889
rect 13 5783 47 5817
rect 85 5783 119 5817
rect 157 5783 191 5817
rect 13 5711 47 5745
rect 85 5711 119 5745
rect 157 5711 191 5745
rect 13 5639 47 5673
rect 85 5639 119 5673
rect 157 5639 191 5673
rect 13 5567 47 5601
rect 85 5567 119 5601
rect 157 5567 191 5601
rect 13 5495 47 5529
rect 85 5495 119 5529
rect 157 5495 191 5529
rect 13 5423 47 5457
rect 85 5423 119 5457
rect 157 5423 191 5457
rect 13 5351 47 5385
rect 85 5351 119 5385
rect 157 5351 191 5385
rect 13 5279 47 5313
rect 85 5279 119 5313
rect 157 5279 191 5313
rect 13 5207 47 5241
rect 85 5207 119 5241
rect 157 5207 191 5241
rect 13 5135 47 5169
rect 85 5135 119 5169
rect 157 5135 191 5169
rect 13 5063 47 5097
rect 85 5063 119 5097
rect 157 5063 191 5097
rect 13 4991 47 5025
rect 85 4991 119 5025
rect 157 4991 191 5025
rect 13 4919 47 4953
rect 85 4919 119 4953
rect 157 4919 191 4953
rect 13 4847 47 4881
rect 85 4847 119 4881
rect 157 4847 191 4881
rect 13 4775 47 4809
rect 85 4775 119 4809
rect 157 4775 191 4809
rect 13 4703 47 4737
rect 85 4703 119 4737
rect 157 4703 191 4737
rect 13 4631 47 4665
rect 85 4631 119 4665
rect 157 4631 191 4665
rect 13 4559 47 4593
rect 85 4559 119 4593
rect 157 4559 191 4593
rect 13 4487 47 4521
rect 85 4487 119 4521
rect 157 4487 191 4521
rect 13 4415 47 4449
rect 85 4415 119 4449
rect 157 4415 191 4449
rect 13 4343 47 4377
rect 85 4343 119 4377
rect 157 4343 191 4377
rect 13 4271 47 4305
rect 85 4271 119 4305
rect 157 4271 191 4305
rect 13 4199 47 4233
rect 85 4199 119 4233
rect 157 4199 191 4233
rect 13 4127 47 4161
rect 85 4127 119 4161
rect 157 4127 191 4161
rect 13 4055 47 4089
rect 85 4055 119 4089
rect 157 4055 191 4089
rect 13 3983 47 4017
rect 85 3983 119 4017
rect 157 3983 191 4017
rect 13 3911 47 3945
rect 85 3911 119 3945
rect 157 3911 191 3945
rect 13 3839 47 3873
rect 85 3839 119 3873
rect 157 3839 191 3873
rect 13 3767 47 3801
rect 85 3767 119 3801
rect 157 3767 191 3801
rect 13 3695 47 3729
rect 85 3695 119 3729
rect 157 3695 191 3729
rect 13 3623 47 3657
rect 85 3623 119 3657
rect 157 3623 191 3657
rect 13 3551 47 3585
rect 85 3551 119 3585
rect 157 3551 191 3585
rect 13 3479 47 3513
rect 85 3479 119 3513
rect 157 3479 191 3513
rect 13 3407 47 3441
rect 85 3407 119 3441
rect 157 3407 191 3441
rect 13 3335 47 3369
rect 85 3335 119 3369
rect 157 3335 191 3369
rect 13 3263 47 3297
rect 85 3263 119 3297
rect 157 3263 191 3297
rect 13 3191 47 3225
rect 85 3191 119 3225
rect 157 3191 191 3225
rect 13 3119 47 3153
rect 85 3119 119 3153
rect 157 3119 191 3153
rect 13 3047 47 3081
rect 85 3047 119 3081
rect 157 3047 191 3081
rect 13 2975 47 3009
rect 85 2975 119 3009
rect 157 2975 191 3009
rect 13 2903 47 2937
rect 85 2903 119 2937
rect 157 2903 191 2937
rect 13 2831 47 2865
rect 85 2831 119 2865
rect 157 2831 191 2865
rect 13 2759 47 2793
rect 85 2759 119 2793
rect 157 2759 191 2793
rect 13 2687 47 2721
rect 85 2687 119 2721
rect 157 2687 191 2721
rect 13 2615 47 2649
rect 85 2615 119 2649
rect 157 2615 191 2649
rect 13 2543 47 2577
rect 85 2543 119 2577
rect 157 2543 191 2577
rect 13 2471 47 2505
rect 85 2471 119 2505
rect 157 2471 191 2505
rect 13 2399 47 2433
rect 85 2399 119 2433
rect 157 2399 191 2433
rect 13 2327 47 2361
rect 85 2327 119 2361
rect 157 2327 191 2361
rect 13 2255 47 2289
rect 85 2255 119 2289
rect 157 2255 191 2289
rect 13 2183 47 2217
rect 85 2183 119 2217
rect 157 2183 191 2217
rect 13 2111 47 2145
rect 85 2111 119 2145
rect 157 2111 191 2145
rect 13 2039 47 2073
rect 85 2039 119 2073
rect 157 2039 191 2073
rect 13 1967 47 2001
rect 85 1967 119 2001
rect 157 1967 191 2001
rect 13 1895 47 1929
rect 85 1895 119 1929
rect 157 1895 191 1929
rect 13 1823 47 1857
rect 85 1823 119 1857
rect 157 1823 191 1857
rect 13 1751 47 1785
rect 85 1751 119 1785
rect 157 1751 191 1785
rect 13 1679 47 1713
rect 85 1679 119 1713
rect 157 1679 191 1713
rect 13 1607 47 1641
rect 85 1607 119 1641
rect 157 1607 191 1641
rect 13 1535 47 1569
rect 85 1535 119 1569
rect 157 1535 191 1569
rect 13 1463 47 1497
rect 85 1463 119 1497
rect 157 1463 191 1497
rect 13 1391 47 1425
rect 85 1391 119 1425
rect 157 1391 191 1425
rect 13 1319 47 1353
rect 85 1319 119 1353
rect 157 1319 191 1353
rect 13 1247 47 1281
rect 85 1247 119 1281
rect 157 1247 191 1281
rect 13 1175 47 1209
rect 85 1175 119 1209
rect 157 1175 191 1209
rect 13 1103 47 1137
rect 85 1103 119 1137
rect 157 1103 191 1137
rect 13 1031 47 1065
rect 85 1031 119 1065
rect 157 1031 191 1065
rect 13 959 47 993
rect 85 959 119 993
rect 157 959 191 993
rect 13 887 47 921
rect 85 887 119 921
rect 157 887 191 921
rect 13 815 47 849
rect 85 815 119 849
rect 157 815 191 849
rect 13 743 47 777
rect 85 743 119 777
rect 157 743 191 777
rect 13 671 47 705
rect 85 671 119 705
rect 157 671 191 705
rect 13 599 47 633
rect 85 599 119 633
rect 157 599 191 633
rect 13 527 47 561
rect 85 527 119 561
rect 157 527 191 561
rect 13 455 47 489
rect 85 455 119 489
rect 157 455 191 489
rect 13 383 47 417
rect 85 383 119 417
rect 157 383 191 417
rect 13 311 47 345
rect 85 311 119 345
rect 157 311 191 345
rect 13 239 47 273
rect 85 239 119 273
rect 157 239 191 273
rect 13 167 47 201
rect 85 167 119 201
rect 157 167 191 201
rect 13 95 47 129
rect 85 95 119 129
rect 157 95 191 129
rect 13 23 47 57
rect 85 23 119 57
rect 157 23 191 57
rect 1017 7943 1051 7977
rect 1089 7943 1123 7977
rect 1161 7943 1195 7977
rect 1017 7871 1051 7905
rect 1089 7871 1123 7905
rect 1161 7871 1195 7905
rect 1017 7799 1051 7833
rect 1089 7799 1123 7833
rect 1161 7799 1195 7833
rect 1017 7727 1051 7761
rect 1089 7727 1123 7761
rect 1161 7727 1195 7761
rect 1017 7655 1051 7689
rect 1089 7655 1123 7689
rect 1161 7655 1195 7689
rect 1017 7583 1051 7617
rect 1089 7583 1123 7617
rect 1161 7583 1195 7617
rect 1017 7511 1051 7545
rect 1089 7511 1123 7545
rect 1161 7511 1195 7545
rect 1017 7439 1051 7473
rect 1089 7439 1123 7473
rect 1161 7439 1195 7473
rect 1017 7367 1051 7401
rect 1089 7367 1123 7401
rect 1161 7367 1195 7401
rect 1017 7295 1051 7329
rect 1089 7295 1123 7329
rect 1161 7295 1195 7329
rect 1017 7223 1051 7257
rect 1089 7223 1123 7257
rect 1161 7223 1195 7257
rect 1017 7151 1051 7185
rect 1089 7151 1123 7185
rect 1161 7151 1195 7185
rect 1017 7079 1051 7113
rect 1089 7079 1123 7113
rect 1161 7079 1195 7113
rect 1017 7007 1051 7041
rect 1089 7007 1123 7041
rect 1161 7007 1195 7041
rect 1017 6935 1051 6969
rect 1089 6935 1123 6969
rect 1161 6935 1195 6969
rect 1017 6863 1051 6897
rect 1089 6863 1123 6897
rect 1161 6863 1195 6897
rect 1017 6791 1051 6825
rect 1089 6791 1123 6825
rect 1161 6791 1195 6825
rect 1017 6719 1051 6753
rect 1089 6719 1123 6753
rect 1161 6719 1195 6753
rect 1017 6647 1051 6681
rect 1089 6647 1123 6681
rect 1161 6647 1195 6681
rect 1017 6575 1051 6609
rect 1089 6575 1123 6609
rect 1161 6575 1195 6609
rect 1017 6503 1051 6537
rect 1089 6503 1123 6537
rect 1161 6503 1195 6537
rect 1017 6431 1051 6465
rect 1089 6431 1123 6465
rect 1161 6431 1195 6465
rect 1017 6359 1051 6393
rect 1089 6359 1123 6393
rect 1161 6359 1195 6393
rect 1017 6287 1051 6321
rect 1089 6287 1123 6321
rect 1161 6287 1195 6321
rect 1017 6215 1051 6249
rect 1089 6215 1123 6249
rect 1161 6215 1195 6249
rect 1017 6143 1051 6177
rect 1089 6143 1123 6177
rect 1161 6143 1195 6177
rect 1017 6071 1051 6105
rect 1089 6071 1123 6105
rect 1161 6071 1195 6105
rect 1017 5999 1051 6033
rect 1089 5999 1123 6033
rect 1161 5999 1195 6033
rect 1017 5927 1051 5961
rect 1089 5927 1123 5961
rect 1161 5927 1195 5961
rect 1017 5855 1051 5889
rect 1089 5855 1123 5889
rect 1161 5855 1195 5889
rect 1017 5783 1051 5817
rect 1089 5783 1123 5817
rect 1161 5783 1195 5817
rect 1017 5711 1051 5745
rect 1089 5711 1123 5745
rect 1161 5711 1195 5745
rect 1017 5639 1051 5673
rect 1089 5639 1123 5673
rect 1161 5639 1195 5673
rect 1017 5567 1051 5601
rect 1089 5567 1123 5601
rect 1161 5567 1195 5601
rect 1017 5495 1051 5529
rect 1089 5495 1123 5529
rect 1161 5495 1195 5529
rect 1017 5423 1051 5457
rect 1089 5423 1123 5457
rect 1161 5423 1195 5457
rect 1017 5351 1051 5385
rect 1089 5351 1123 5385
rect 1161 5351 1195 5385
rect 1017 5279 1051 5313
rect 1089 5279 1123 5313
rect 1161 5279 1195 5313
rect 1017 5207 1051 5241
rect 1089 5207 1123 5241
rect 1161 5207 1195 5241
rect 1017 5135 1051 5169
rect 1089 5135 1123 5169
rect 1161 5135 1195 5169
rect 1017 5063 1051 5097
rect 1089 5063 1123 5097
rect 1161 5063 1195 5097
rect 1017 4991 1051 5025
rect 1089 4991 1123 5025
rect 1161 4991 1195 5025
rect 1017 4919 1051 4953
rect 1089 4919 1123 4953
rect 1161 4919 1195 4953
rect 1017 4847 1051 4881
rect 1089 4847 1123 4881
rect 1161 4847 1195 4881
rect 1017 4775 1051 4809
rect 1089 4775 1123 4809
rect 1161 4775 1195 4809
rect 1017 4703 1051 4737
rect 1089 4703 1123 4737
rect 1161 4703 1195 4737
rect 1017 4631 1051 4665
rect 1089 4631 1123 4665
rect 1161 4631 1195 4665
rect 1017 4559 1051 4593
rect 1089 4559 1123 4593
rect 1161 4559 1195 4593
rect 1017 4487 1051 4521
rect 1089 4487 1123 4521
rect 1161 4487 1195 4521
rect 1017 4415 1051 4449
rect 1089 4415 1123 4449
rect 1161 4415 1195 4449
rect 1017 4343 1051 4377
rect 1089 4343 1123 4377
rect 1161 4343 1195 4377
rect 1017 4271 1051 4305
rect 1089 4271 1123 4305
rect 1161 4271 1195 4305
rect 1017 4199 1051 4233
rect 1089 4199 1123 4233
rect 1161 4199 1195 4233
rect 1017 4127 1051 4161
rect 1089 4127 1123 4161
rect 1161 4127 1195 4161
rect 1017 4055 1051 4089
rect 1089 4055 1123 4089
rect 1161 4055 1195 4089
rect 1017 3983 1051 4017
rect 1089 3983 1123 4017
rect 1161 3983 1195 4017
rect 1017 3911 1051 3945
rect 1089 3911 1123 3945
rect 1161 3911 1195 3945
rect 1017 3839 1051 3873
rect 1089 3839 1123 3873
rect 1161 3839 1195 3873
rect 1017 3767 1051 3801
rect 1089 3767 1123 3801
rect 1161 3767 1195 3801
rect 1017 3695 1051 3729
rect 1089 3695 1123 3729
rect 1161 3695 1195 3729
rect 1017 3623 1051 3657
rect 1089 3623 1123 3657
rect 1161 3623 1195 3657
rect 1017 3551 1051 3585
rect 1089 3551 1123 3585
rect 1161 3551 1195 3585
rect 1017 3479 1051 3513
rect 1089 3479 1123 3513
rect 1161 3479 1195 3513
rect 1017 3407 1051 3441
rect 1089 3407 1123 3441
rect 1161 3407 1195 3441
rect 1017 3335 1051 3369
rect 1089 3335 1123 3369
rect 1161 3335 1195 3369
rect 1017 3263 1051 3297
rect 1089 3263 1123 3297
rect 1161 3263 1195 3297
rect 1017 3191 1051 3225
rect 1089 3191 1123 3225
rect 1161 3191 1195 3225
rect 1017 3119 1051 3153
rect 1089 3119 1123 3153
rect 1161 3119 1195 3153
rect 1017 3047 1051 3081
rect 1089 3047 1123 3081
rect 1161 3047 1195 3081
rect 1017 2975 1051 3009
rect 1089 2975 1123 3009
rect 1161 2975 1195 3009
rect 1017 2903 1051 2937
rect 1089 2903 1123 2937
rect 1161 2903 1195 2937
rect 1017 2831 1051 2865
rect 1089 2831 1123 2865
rect 1161 2831 1195 2865
rect 1017 2759 1051 2793
rect 1089 2759 1123 2793
rect 1161 2759 1195 2793
rect 1017 2687 1051 2721
rect 1089 2687 1123 2721
rect 1161 2687 1195 2721
rect 1017 2615 1051 2649
rect 1089 2615 1123 2649
rect 1161 2615 1195 2649
rect 1017 2543 1051 2577
rect 1089 2543 1123 2577
rect 1161 2543 1195 2577
rect 1017 2471 1051 2505
rect 1089 2471 1123 2505
rect 1161 2471 1195 2505
rect 1017 2399 1051 2433
rect 1089 2399 1123 2433
rect 1161 2399 1195 2433
rect 1017 2327 1051 2361
rect 1089 2327 1123 2361
rect 1161 2327 1195 2361
rect 1017 2255 1051 2289
rect 1089 2255 1123 2289
rect 1161 2255 1195 2289
rect 1017 2183 1051 2217
rect 1089 2183 1123 2217
rect 1161 2183 1195 2217
rect 1017 2111 1051 2145
rect 1089 2111 1123 2145
rect 1161 2111 1195 2145
rect 1017 2039 1051 2073
rect 1089 2039 1123 2073
rect 1161 2039 1195 2073
rect 1017 1967 1051 2001
rect 1089 1967 1123 2001
rect 1161 1967 1195 2001
rect 1017 1895 1051 1929
rect 1089 1895 1123 1929
rect 1161 1895 1195 1929
rect 1017 1823 1051 1857
rect 1089 1823 1123 1857
rect 1161 1823 1195 1857
rect 1017 1751 1051 1785
rect 1089 1751 1123 1785
rect 1161 1751 1195 1785
rect 1017 1679 1051 1713
rect 1089 1679 1123 1713
rect 1161 1679 1195 1713
rect 1017 1607 1051 1641
rect 1089 1607 1123 1641
rect 1161 1607 1195 1641
rect 1017 1535 1051 1569
rect 1089 1535 1123 1569
rect 1161 1535 1195 1569
rect 1017 1463 1051 1497
rect 1089 1463 1123 1497
rect 1161 1463 1195 1497
rect 1017 1391 1051 1425
rect 1089 1391 1123 1425
rect 1161 1391 1195 1425
rect 1017 1319 1051 1353
rect 1089 1319 1123 1353
rect 1161 1319 1195 1353
rect 1017 1247 1051 1281
rect 1089 1247 1123 1281
rect 1161 1247 1195 1281
rect 1017 1175 1051 1209
rect 1089 1175 1123 1209
rect 1161 1175 1195 1209
rect 1017 1103 1051 1137
rect 1089 1103 1123 1137
rect 1161 1103 1195 1137
rect 1017 1031 1051 1065
rect 1089 1031 1123 1065
rect 1161 1031 1195 1065
rect 1017 959 1051 993
rect 1089 959 1123 993
rect 1161 959 1195 993
rect 1017 887 1051 921
rect 1089 887 1123 921
rect 1161 887 1195 921
rect 1017 815 1051 849
rect 1089 815 1123 849
rect 1161 815 1195 849
rect 1017 743 1051 777
rect 1089 743 1123 777
rect 1161 743 1195 777
rect 1017 671 1051 705
rect 1089 671 1123 705
rect 1161 671 1195 705
rect 1017 599 1051 633
rect 1089 599 1123 633
rect 1161 599 1195 633
rect 1017 527 1051 561
rect 1089 527 1123 561
rect 1161 527 1195 561
rect 1017 455 1051 489
rect 1089 455 1123 489
rect 1161 455 1195 489
rect 1017 383 1051 417
rect 1089 383 1123 417
rect 1161 383 1195 417
rect 1017 311 1051 345
rect 1089 311 1123 345
rect 1161 311 1195 345
rect 1017 239 1051 273
rect 1089 239 1123 273
rect 1161 239 1195 273
rect 1017 167 1051 201
rect 1089 167 1123 201
rect 1161 167 1195 201
rect 1017 95 1051 129
rect 1089 95 1123 129
rect 1161 95 1195 129
rect 1017 23 1051 57
rect 1089 23 1123 57
rect 1161 23 1195 57
<< nsubdiff >>
rect 1208 7977 1473 8000
rect 1208 7943 1252 7977
rect 1286 7943 1324 7977
rect 1358 7943 1396 7977
rect 1430 7943 1473 7977
rect 1208 7905 1473 7943
rect 1208 7871 1252 7905
rect 1286 7871 1324 7905
rect 1358 7871 1396 7905
rect 1430 7871 1473 7905
rect 1208 7833 1473 7871
rect 1208 7799 1252 7833
rect 1286 7799 1324 7833
rect 1358 7799 1396 7833
rect 1430 7799 1473 7833
rect 1208 7761 1473 7799
rect 1208 7727 1252 7761
rect 1286 7727 1324 7761
rect 1358 7727 1396 7761
rect 1430 7727 1473 7761
rect 1208 7689 1473 7727
rect 1208 7655 1252 7689
rect 1286 7655 1324 7689
rect 1358 7655 1396 7689
rect 1430 7655 1473 7689
rect 1208 7617 1473 7655
rect 1208 7583 1252 7617
rect 1286 7583 1324 7617
rect 1358 7583 1396 7617
rect 1430 7583 1473 7617
rect 1208 7545 1473 7583
rect 1208 7511 1252 7545
rect 1286 7511 1324 7545
rect 1358 7511 1396 7545
rect 1430 7511 1473 7545
rect 1208 7473 1473 7511
rect 1208 7439 1252 7473
rect 1286 7439 1324 7473
rect 1358 7439 1396 7473
rect 1430 7439 1473 7473
rect 1208 7401 1473 7439
rect 1208 7367 1252 7401
rect 1286 7367 1324 7401
rect 1358 7367 1396 7401
rect 1430 7367 1473 7401
rect 1208 7329 1473 7367
rect 1208 7295 1252 7329
rect 1286 7295 1324 7329
rect 1358 7295 1396 7329
rect 1430 7295 1473 7329
rect 1208 7257 1473 7295
rect 1208 7223 1252 7257
rect 1286 7223 1324 7257
rect 1358 7223 1396 7257
rect 1430 7223 1473 7257
rect 1208 7185 1473 7223
rect 1208 7151 1252 7185
rect 1286 7151 1324 7185
rect 1358 7151 1396 7185
rect 1430 7151 1473 7185
rect 1208 7113 1473 7151
rect 1208 7079 1252 7113
rect 1286 7079 1324 7113
rect 1358 7079 1396 7113
rect 1430 7079 1473 7113
rect 1208 7041 1473 7079
rect 1208 7007 1252 7041
rect 1286 7007 1324 7041
rect 1358 7007 1396 7041
rect 1430 7007 1473 7041
rect 1208 6969 1473 7007
rect 1208 6935 1252 6969
rect 1286 6935 1324 6969
rect 1358 6935 1396 6969
rect 1430 6935 1473 6969
rect 1208 6897 1473 6935
rect 1208 6863 1252 6897
rect 1286 6863 1324 6897
rect 1358 6863 1396 6897
rect 1430 6863 1473 6897
rect 1208 6825 1473 6863
rect 1208 6791 1252 6825
rect 1286 6791 1324 6825
rect 1358 6791 1396 6825
rect 1430 6791 1473 6825
rect 1208 6753 1473 6791
rect 1208 6719 1252 6753
rect 1286 6719 1324 6753
rect 1358 6719 1396 6753
rect 1430 6719 1473 6753
rect 1208 6681 1473 6719
rect 1208 6647 1252 6681
rect 1286 6647 1324 6681
rect 1358 6647 1396 6681
rect 1430 6647 1473 6681
rect 1208 6609 1473 6647
rect 1208 6575 1252 6609
rect 1286 6575 1324 6609
rect 1358 6575 1396 6609
rect 1430 6575 1473 6609
rect 1208 6537 1473 6575
rect 1208 6503 1252 6537
rect 1286 6503 1324 6537
rect 1358 6503 1396 6537
rect 1430 6503 1473 6537
rect 1208 6465 1473 6503
rect 1208 6431 1252 6465
rect 1286 6431 1324 6465
rect 1358 6431 1396 6465
rect 1430 6431 1473 6465
rect 1208 6393 1473 6431
rect 1208 6359 1252 6393
rect 1286 6359 1324 6393
rect 1358 6359 1396 6393
rect 1430 6359 1473 6393
rect 1208 6321 1473 6359
rect 1208 6287 1252 6321
rect 1286 6287 1324 6321
rect 1358 6287 1396 6321
rect 1430 6287 1473 6321
rect 1208 6249 1473 6287
rect 1208 6215 1252 6249
rect 1286 6215 1324 6249
rect 1358 6215 1396 6249
rect 1430 6215 1473 6249
rect 1208 6177 1473 6215
rect 1208 6143 1252 6177
rect 1286 6143 1324 6177
rect 1358 6143 1396 6177
rect 1430 6143 1473 6177
rect 1208 6105 1473 6143
rect 1208 6071 1252 6105
rect 1286 6071 1324 6105
rect 1358 6071 1396 6105
rect 1430 6071 1473 6105
rect 1208 6033 1473 6071
rect 1208 5999 1252 6033
rect 1286 5999 1324 6033
rect 1358 5999 1396 6033
rect 1430 5999 1473 6033
rect 1208 5961 1473 5999
rect 1208 5927 1252 5961
rect 1286 5927 1324 5961
rect 1358 5927 1396 5961
rect 1430 5927 1473 5961
rect 1208 5889 1473 5927
rect 1208 5855 1252 5889
rect 1286 5855 1324 5889
rect 1358 5855 1396 5889
rect 1430 5855 1473 5889
rect 1208 5817 1473 5855
rect 1208 5783 1252 5817
rect 1286 5783 1324 5817
rect 1358 5783 1396 5817
rect 1430 5783 1473 5817
rect 1208 5745 1473 5783
rect 1208 5711 1252 5745
rect 1286 5711 1324 5745
rect 1358 5711 1396 5745
rect 1430 5711 1473 5745
rect 1208 5673 1473 5711
rect 1208 5639 1252 5673
rect 1286 5639 1324 5673
rect 1358 5639 1396 5673
rect 1430 5639 1473 5673
rect 1208 5601 1473 5639
rect 1208 5567 1252 5601
rect 1286 5567 1324 5601
rect 1358 5567 1396 5601
rect 1430 5567 1473 5601
rect 1208 5529 1473 5567
rect 1208 5495 1252 5529
rect 1286 5495 1324 5529
rect 1358 5495 1396 5529
rect 1430 5495 1473 5529
rect 1208 5457 1473 5495
rect 1208 5423 1252 5457
rect 1286 5423 1324 5457
rect 1358 5423 1396 5457
rect 1430 5423 1473 5457
rect 1208 5385 1473 5423
rect 1208 5351 1252 5385
rect 1286 5351 1324 5385
rect 1358 5351 1396 5385
rect 1430 5351 1473 5385
rect 1208 5313 1473 5351
rect 1208 5279 1252 5313
rect 1286 5279 1324 5313
rect 1358 5279 1396 5313
rect 1430 5279 1473 5313
rect 1208 5241 1473 5279
rect 1208 5207 1252 5241
rect 1286 5207 1324 5241
rect 1358 5207 1396 5241
rect 1430 5207 1473 5241
rect 1208 5169 1473 5207
rect 1208 5135 1252 5169
rect 1286 5135 1324 5169
rect 1358 5135 1396 5169
rect 1430 5135 1473 5169
rect 1208 5097 1473 5135
rect 1208 5063 1252 5097
rect 1286 5063 1324 5097
rect 1358 5063 1396 5097
rect 1430 5063 1473 5097
rect 1208 5025 1473 5063
rect 1208 4991 1252 5025
rect 1286 4991 1324 5025
rect 1358 4991 1396 5025
rect 1430 4991 1473 5025
rect 1208 4953 1473 4991
rect 1208 4919 1252 4953
rect 1286 4919 1324 4953
rect 1358 4919 1396 4953
rect 1430 4919 1473 4953
rect 1208 4881 1473 4919
rect 1208 4847 1252 4881
rect 1286 4847 1324 4881
rect 1358 4847 1396 4881
rect 1430 4847 1473 4881
rect 1208 4809 1473 4847
rect 1208 4775 1252 4809
rect 1286 4775 1324 4809
rect 1358 4775 1396 4809
rect 1430 4775 1473 4809
rect 1208 4737 1473 4775
rect 1208 4703 1252 4737
rect 1286 4703 1324 4737
rect 1358 4703 1396 4737
rect 1430 4703 1473 4737
rect 1208 4665 1473 4703
rect 1208 4631 1252 4665
rect 1286 4631 1324 4665
rect 1358 4631 1396 4665
rect 1430 4631 1473 4665
rect 1208 4593 1473 4631
rect 1208 4559 1252 4593
rect 1286 4559 1324 4593
rect 1358 4559 1396 4593
rect 1430 4559 1473 4593
rect 1208 4521 1473 4559
rect 1208 4487 1252 4521
rect 1286 4487 1324 4521
rect 1358 4487 1396 4521
rect 1430 4487 1473 4521
rect 1208 4449 1473 4487
rect 1208 4415 1252 4449
rect 1286 4415 1324 4449
rect 1358 4415 1396 4449
rect 1430 4415 1473 4449
rect 1208 4377 1473 4415
rect 1208 4343 1252 4377
rect 1286 4343 1324 4377
rect 1358 4343 1396 4377
rect 1430 4343 1473 4377
rect 1208 4305 1473 4343
rect 1208 4271 1252 4305
rect 1286 4271 1324 4305
rect 1358 4271 1396 4305
rect 1430 4271 1473 4305
rect 1208 4233 1473 4271
rect 1208 4199 1252 4233
rect 1286 4199 1324 4233
rect 1358 4199 1396 4233
rect 1430 4199 1473 4233
rect 1208 4161 1473 4199
rect 1208 4127 1252 4161
rect 1286 4127 1324 4161
rect 1358 4127 1396 4161
rect 1430 4127 1473 4161
rect 1208 4089 1473 4127
rect 1208 4055 1252 4089
rect 1286 4055 1324 4089
rect 1358 4055 1396 4089
rect 1430 4055 1473 4089
rect 1208 4017 1473 4055
rect 1208 3983 1252 4017
rect 1286 3983 1324 4017
rect 1358 3983 1396 4017
rect 1430 3983 1473 4017
rect 1208 3945 1473 3983
rect 1208 3911 1252 3945
rect 1286 3911 1324 3945
rect 1358 3911 1396 3945
rect 1430 3911 1473 3945
rect 1208 3873 1473 3911
rect 1208 3839 1252 3873
rect 1286 3839 1324 3873
rect 1358 3839 1396 3873
rect 1430 3839 1473 3873
rect 1208 3801 1473 3839
rect 1208 3767 1252 3801
rect 1286 3767 1324 3801
rect 1358 3767 1396 3801
rect 1430 3767 1473 3801
rect 1208 3729 1473 3767
rect 1208 3695 1252 3729
rect 1286 3695 1324 3729
rect 1358 3695 1396 3729
rect 1430 3695 1473 3729
rect 1208 3657 1473 3695
rect 1208 3623 1252 3657
rect 1286 3623 1324 3657
rect 1358 3623 1396 3657
rect 1430 3623 1473 3657
rect 1208 3585 1473 3623
rect 1208 3551 1252 3585
rect 1286 3551 1324 3585
rect 1358 3551 1396 3585
rect 1430 3551 1473 3585
rect 1208 3513 1473 3551
rect 1208 3479 1252 3513
rect 1286 3479 1324 3513
rect 1358 3479 1396 3513
rect 1430 3479 1473 3513
rect 1208 3441 1473 3479
rect 1208 3407 1252 3441
rect 1286 3407 1324 3441
rect 1358 3407 1396 3441
rect 1430 3407 1473 3441
rect 1208 3369 1473 3407
rect 1208 3335 1252 3369
rect 1286 3335 1324 3369
rect 1358 3335 1396 3369
rect 1430 3335 1473 3369
rect 1208 3297 1473 3335
rect 1208 3263 1252 3297
rect 1286 3263 1324 3297
rect 1358 3263 1396 3297
rect 1430 3263 1473 3297
rect 1208 3225 1473 3263
rect 1208 3191 1252 3225
rect 1286 3191 1324 3225
rect 1358 3191 1396 3225
rect 1430 3191 1473 3225
rect 1208 3153 1473 3191
rect 1208 3119 1252 3153
rect 1286 3119 1324 3153
rect 1358 3119 1396 3153
rect 1430 3119 1473 3153
rect 1208 3081 1473 3119
rect 1208 3047 1252 3081
rect 1286 3047 1324 3081
rect 1358 3047 1396 3081
rect 1430 3047 1473 3081
rect 1208 3009 1473 3047
rect 1208 2975 1252 3009
rect 1286 2975 1324 3009
rect 1358 2975 1396 3009
rect 1430 2975 1473 3009
rect 1208 2937 1473 2975
rect 1208 2903 1252 2937
rect 1286 2903 1324 2937
rect 1358 2903 1396 2937
rect 1430 2903 1473 2937
rect 1208 2865 1473 2903
rect 1208 2831 1252 2865
rect 1286 2831 1324 2865
rect 1358 2831 1396 2865
rect 1430 2831 1473 2865
rect 1208 2793 1473 2831
rect 1208 2759 1252 2793
rect 1286 2759 1324 2793
rect 1358 2759 1396 2793
rect 1430 2759 1473 2793
rect 1208 2721 1473 2759
rect 1208 2687 1252 2721
rect 1286 2687 1324 2721
rect 1358 2687 1396 2721
rect 1430 2687 1473 2721
rect 1208 2649 1473 2687
rect 1208 2615 1252 2649
rect 1286 2615 1324 2649
rect 1358 2615 1396 2649
rect 1430 2615 1473 2649
rect 1208 2577 1473 2615
rect 1208 2543 1252 2577
rect 1286 2543 1324 2577
rect 1358 2543 1396 2577
rect 1430 2543 1473 2577
rect 1208 2505 1473 2543
rect 1208 2471 1252 2505
rect 1286 2471 1324 2505
rect 1358 2471 1396 2505
rect 1430 2471 1473 2505
rect 1208 2433 1473 2471
rect 1208 2399 1252 2433
rect 1286 2399 1324 2433
rect 1358 2399 1396 2433
rect 1430 2399 1473 2433
rect 1208 2361 1473 2399
rect 1208 2327 1252 2361
rect 1286 2327 1324 2361
rect 1358 2327 1396 2361
rect 1430 2327 1473 2361
rect 1208 2289 1473 2327
rect 1208 2255 1252 2289
rect 1286 2255 1324 2289
rect 1358 2255 1396 2289
rect 1430 2255 1473 2289
rect 1208 2217 1473 2255
rect 1208 2183 1252 2217
rect 1286 2183 1324 2217
rect 1358 2183 1396 2217
rect 1430 2183 1473 2217
rect 1208 2145 1473 2183
rect 1208 2111 1252 2145
rect 1286 2111 1324 2145
rect 1358 2111 1396 2145
rect 1430 2111 1473 2145
rect 1208 2073 1473 2111
rect 1208 2039 1252 2073
rect 1286 2039 1324 2073
rect 1358 2039 1396 2073
rect 1430 2039 1473 2073
rect 1208 2001 1473 2039
rect 1208 1967 1252 2001
rect 1286 1967 1324 2001
rect 1358 1967 1396 2001
rect 1430 1967 1473 2001
rect 1208 1929 1473 1967
rect 1208 1895 1252 1929
rect 1286 1895 1324 1929
rect 1358 1895 1396 1929
rect 1430 1895 1473 1929
rect 1208 1857 1473 1895
rect 1208 1823 1252 1857
rect 1286 1823 1324 1857
rect 1358 1823 1396 1857
rect 1430 1823 1473 1857
rect 1208 1785 1473 1823
rect 1208 1751 1252 1785
rect 1286 1751 1324 1785
rect 1358 1751 1396 1785
rect 1430 1751 1473 1785
rect 1208 1713 1473 1751
rect 1208 1679 1252 1713
rect 1286 1679 1324 1713
rect 1358 1679 1396 1713
rect 1430 1679 1473 1713
rect 1208 1641 1473 1679
rect 1208 1607 1252 1641
rect 1286 1607 1324 1641
rect 1358 1607 1396 1641
rect 1430 1607 1473 1641
rect 1208 1569 1473 1607
rect 1208 1535 1252 1569
rect 1286 1535 1324 1569
rect 1358 1535 1396 1569
rect 1430 1535 1473 1569
rect 1208 1497 1473 1535
rect 1208 1463 1252 1497
rect 1286 1463 1324 1497
rect 1358 1463 1396 1497
rect 1430 1463 1473 1497
rect 1208 1425 1473 1463
rect 1208 1391 1252 1425
rect 1286 1391 1324 1425
rect 1358 1391 1396 1425
rect 1430 1391 1473 1425
rect 1208 1353 1473 1391
rect 1208 1319 1252 1353
rect 1286 1319 1324 1353
rect 1358 1319 1396 1353
rect 1430 1319 1473 1353
rect 1208 1281 1473 1319
rect 1208 1247 1252 1281
rect 1286 1247 1324 1281
rect 1358 1247 1396 1281
rect 1430 1247 1473 1281
rect 1208 1209 1473 1247
rect 1208 1175 1252 1209
rect 1286 1175 1324 1209
rect 1358 1175 1396 1209
rect 1430 1175 1473 1209
rect 1208 1137 1473 1175
rect 1208 1103 1252 1137
rect 1286 1103 1324 1137
rect 1358 1103 1396 1137
rect 1430 1103 1473 1137
rect 1208 1065 1473 1103
rect 1208 1031 1252 1065
rect 1286 1031 1324 1065
rect 1358 1031 1396 1065
rect 1430 1031 1473 1065
rect 1208 993 1473 1031
rect 1208 959 1252 993
rect 1286 959 1324 993
rect 1358 959 1396 993
rect 1430 959 1473 993
rect 1208 921 1473 959
rect 1208 887 1252 921
rect 1286 887 1324 921
rect 1358 887 1396 921
rect 1430 887 1473 921
rect 1208 849 1473 887
rect 1208 815 1252 849
rect 1286 815 1324 849
rect 1358 815 1396 849
rect 1430 815 1473 849
rect 1208 777 1473 815
rect 1208 743 1252 777
rect 1286 743 1324 777
rect 1358 743 1396 777
rect 1430 743 1473 777
rect 1208 705 1473 743
rect 1208 671 1252 705
rect 1286 671 1324 705
rect 1358 671 1396 705
rect 1430 671 1473 705
rect 1208 633 1473 671
rect 1208 599 1252 633
rect 1286 599 1324 633
rect 1358 599 1396 633
rect 1430 599 1473 633
rect 1208 561 1473 599
rect 1208 527 1252 561
rect 1286 527 1324 561
rect 1358 527 1396 561
rect 1430 527 1473 561
rect 1208 489 1473 527
rect 1208 455 1252 489
rect 1286 455 1324 489
rect 1358 455 1396 489
rect 1430 455 1473 489
rect 1208 417 1473 455
rect 1208 383 1252 417
rect 1286 383 1324 417
rect 1358 383 1396 417
rect 1430 383 1473 417
rect 1208 345 1473 383
rect 1208 311 1252 345
rect 1286 311 1324 345
rect 1358 311 1396 345
rect 1430 311 1473 345
rect 1208 273 1473 311
rect 1208 239 1252 273
rect 1286 239 1324 273
rect 1358 239 1396 273
rect 1430 239 1473 273
rect 1208 201 1473 239
rect 1208 167 1252 201
rect 1286 167 1324 201
rect 1358 167 1396 201
rect 1430 167 1473 201
rect 1208 129 1473 167
rect 1208 95 1252 129
rect 1286 95 1324 129
rect 1358 95 1396 129
rect 1430 95 1473 129
rect 1208 57 1473 95
rect 1208 23 1252 57
rect 1286 23 1324 57
rect 1358 23 1396 57
rect 1430 23 1473 57
rect 1208 0 1473 23
<< nsubdiffcont >>
rect 1252 7943 1286 7977
rect 1324 7943 1358 7977
rect 1396 7943 1430 7977
rect 1252 7871 1286 7905
rect 1324 7871 1358 7905
rect 1396 7871 1430 7905
rect 1252 7799 1286 7833
rect 1324 7799 1358 7833
rect 1396 7799 1430 7833
rect 1252 7727 1286 7761
rect 1324 7727 1358 7761
rect 1396 7727 1430 7761
rect 1252 7655 1286 7689
rect 1324 7655 1358 7689
rect 1396 7655 1430 7689
rect 1252 7583 1286 7617
rect 1324 7583 1358 7617
rect 1396 7583 1430 7617
rect 1252 7511 1286 7545
rect 1324 7511 1358 7545
rect 1396 7511 1430 7545
rect 1252 7439 1286 7473
rect 1324 7439 1358 7473
rect 1396 7439 1430 7473
rect 1252 7367 1286 7401
rect 1324 7367 1358 7401
rect 1396 7367 1430 7401
rect 1252 7295 1286 7329
rect 1324 7295 1358 7329
rect 1396 7295 1430 7329
rect 1252 7223 1286 7257
rect 1324 7223 1358 7257
rect 1396 7223 1430 7257
rect 1252 7151 1286 7185
rect 1324 7151 1358 7185
rect 1396 7151 1430 7185
rect 1252 7079 1286 7113
rect 1324 7079 1358 7113
rect 1396 7079 1430 7113
rect 1252 7007 1286 7041
rect 1324 7007 1358 7041
rect 1396 7007 1430 7041
rect 1252 6935 1286 6969
rect 1324 6935 1358 6969
rect 1396 6935 1430 6969
rect 1252 6863 1286 6897
rect 1324 6863 1358 6897
rect 1396 6863 1430 6897
rect 1252 6791 1286 6825
rect 1324 6791 1358 6825
rect 1396 6791 1430 6825
rect 1252 6719 1286 6753
rect 1324 6719 1358 6753
rect 1396 6719 1430 6753
rect 1252 6647 1286 6681
rect 1324 6647 1358 6681
rect 1396 6647 1430 6681
rect 1252 6575 1286 6609
rect 1324 6575 1358 6609
rect 1396 6575 1430 6609
rect 1252 6503 1286 6537
rect 1324 6503 1358 6537
rect 1396 6503 1430 6537
rect 1252 6431 1286 6465
rect 1324 6431 1358 6465
rect 1396 6431 1430 6465
rect 1252 6359 1286 6393
rect 1324 6359 1358 6393
rect 1396 6359 1430 6393
rect 1252 6287 1286 6321
rect 1324 6287 1358 6321
rect 1396 6287 1430 6321
rect 1252 6215 1286 6249
rect 1324 6215 1358 6249
rect 1396 6215 1430 6249
rect 1252 6143 1286 6177
rect 1324 6143 1358 6177
rect 1396 6143 1430 6177
rect 1252 6071 1286 6105
rect 1324 6071 1358 6105
rect 1396 6071 1430 6105
rect 1252 5999 1286 6033
rect 1324 5999 1358 6033
rect 1396 5999 1430 6033
rect 1252 5927 1286 5961
rect 1324 5927 1358 5961
rect 1396 5927 1430 5961
rect 1252 5855 1286 5889
rect 1324 5855 1358 5889
rect 1396 5855 1430 5889
rect 1252 5783 1286 5817
rect 1324 5783 1358 5817
rect 1396 5783 1430 5817
rect 1252 5711 1286 5745
rect 1324 5711 1358 5745
rect 1396 5711 1430 5745
rect 1252 5639 1286 5673
rect 1324 5639 1358 5673
rect 1396 5639 1430 5673
rect 1252 5567 1286 5601
rect 1324 5567 1358 5601
rect 1396 5567 1430 5601
rect 1252 5495 1286 5529
rect 1324 5495 1358 5529
rect 1396 5495 1430 5529
rect 1252 5423 1286 5457
rect 1324 5423 1358 5457
rect 1396 5423 1430 5457
rect 1252 5351 1286 5385
rect 1324 5351 1358 5385
rect 1396 5351 1430 5385
rect 1252 5279 1286 5313
rect 1324 5279 1358 5313
rect 1396 5279 1430 5313
rect 1252 5207 1286 5241
rect 1324 5207 1358 5241
rect 1396 5207 1430 5241
rect 1252 5135 1286 5169
rect 1324 5135 1358 5169
rect 1396 5135 1430 5169
rect 1252 5063 1286 5097
rect 1324 5063 1358 5097
rect 1396 5063 1430 5097
rect 1252 4991 1286 5025
rect 1324 4991 1358 5025
rect 1396 4991 1430 5025
rect 1252 4919 1286 4953
rect 1324 4919 1358 4953
rect 1396 4919 1430 4953
rect 1252 4847 1286 4881
rect 1324 4847 1358 4881
rect 1396 4847 1430 4881
rect 1252 4775 1286 4809
rect 1324 4775 1358 4809
rect 1396 4775 1430 4809
rect 1252 4703 1286 4737
rect 1324 4703 1358 4737
rect 1396 4703 1430 4737
rect 1252 4631 1286 4665
rect 1324 4631 1358 4665
rect 1396 4631 1430 4665
rect 1252 4559 1286 4593
rect 1324 4559 1358 4593
rect 1396 4559 1430 4593
rect 1252 4487 1286 4521
rect 1324 4487 1358 4521
rect 1396 4487 1430 4521
rect 1252 4415 1286 4449
rect 1324 4415 1358 4449
rect 1396 4415 1430 4449
rect 1252 4343 1286 4377
rect 1324 4343 1358 4377
rect 1396 4343 1430 4377
rect 1252 4271 1286 4305
rect 1324 4271 1358 4305
rect 1396 4271 1430 4305
rect 1252 4199 1286 4233
rect 1324 4199 1358 4233
rect 1396 4199 1430 4233
rect 1252 4127 1286 4161
rect 1324 4127 1358 4161
rect 1396 4127 1430 4161
rect 1252 4055 1286 4089
rect 1324 4055 1358 4089
rect 1396 4055 1430 4089
rect 1252 3983 1286 4017
rect 1324 3983 1358 4017
rect 1396 3983 1430 4017
rect 1252 3911 1286 3945
rect 1324 3911 1358 3945
rect 1396 3911 1430 3945
rect 1252 3839 1286 3873
rect 1324 3839 1358 3873
rect 1396 3839 1430 3873
rect 1252 3767 1286 3801
rect 1324 3767 1358 3801
rect 1396 3767 1430 3801
rect 1252 3695 1286 3729
rect 1324 3695 1358 3729
rect 1396 3695 1430 3729
rect 1252 3623 1286 3657
rect 1324 3623 1358 3657
rect 1396 3623 1430 3657
rect 1252 3551 1286 3585
rect 1324 3551 1358 3585
rect 1396 3551 1430 3585
rect 1252 3479 1286 3513
rect 1324 3479 1358 3513
rect 1396 3479 1430 3513
rect 1252 3407 1286 3441
rect 1324 3407 1358 3441
rect 1396 3407 1430 3441
rect 1252 3335 1286 3369
rect 1324 3335 1358 3369
rect 1396 3335 1430 3369
rect 1252 3263 1286 3297
rect 1324 3263 1358 3297
rect 1396 3263 1430 3297
rect 1252 3191 1286 3225
rect 1324 3191 1358 3225
rect 1396 3191 1430 3225
rect 1252 3119 1286 3153
rect 1324 3119 1358 3153
rect 1396 3119 1430 3153
rect 1252 3047 1286 3081
rect 1324 3047 1358 3081
rect 1396 3047 1430 3081
rect 1252 2975 1286 3009
rect 1324 2975 1358 3009
rect 1396 2975 1430 3009
rect 1252 2903 1286 2937
rect 1324 2903 1358 2937
rect 1396 2903 1430 2937
rect 1252 2831 1286 2865
rect 1324 2831 1358 2865
rect 1396 2831 1430 2865
rect 1252 2759 1286 2793
rect 1324 2759 1358 2793
rect 1396 2759 1430 2793
rect 1252 2687 1286 2721
rect 1324 2687 1358 2721
rect 1396 2687 1430 2721
rect 1252 2615 1286 2649
rect 1324 2615 1358 2649
rect 1396 2615 1430 2649
rect 1252 2543 1286 2577
rect 1324 2543 1358 2577
rect 1396 2543 1430 2577
rect 1252 2471 1286 2505
rect 1324 2471 1358 2505
rect 1396 2471 1430 2505
rect 1252 2399 1286 2433
rect 1324 2399 1358 2433
rect 1396 2399 1430 2433
rect 1252 2327 1286 2361
rect 1324 2327 1358 2361
rect 1396 2327 1430 2361
rect 1252 2255 1286 2289
rect 1324 2255 1358 2289
rect 1396 2255 1430 2289
rect 1252 2183 1286 2217
rect 1324 2183 1358 2217
rect 1396 2183 1430 2217
rect 1252 2111 1286 2145
rect 1324 2111 1358 2145
rect 1396 2111 1430 2145
rect 1252 2039 1286 2073
rect 1324 2039 1358 2073
rect 1396 2039 1430 2073
rect 1252 1967 1286 2001
rect 1324 1967 1358 2001
rect 1396 1967 1430 2001
rect 1252 1895 1286 1929
rect 1324 1895 1358 1929
rect 1396 1895 1430 1929
rect 1252 1823 1286 1857
rect 1324 1823 1358 1857
rect 1396 1823 1430 1857
rect 1252 1751 1286 1785
rect 1324 1751 1358 1785
rect 1396 1751 1430 1785
rect 1252 1679 1286 1713
rect 1324 1679 1358 1713
rect 1396 1679 1430 1713
rect 1252 1607 1286 1641
rect 1324 1607 1358 1641
rect 1396 1607 1430 1641
rect 1252 1535 1286 1569
rect 1324 1535 1358 1569
rect 1396 1535 1430 1569
rect 1252 1463 1286 1497
rect 1324 1463 1358 1497
rect 1396 1463 1430 1497
rect 1252 1391 1286 1425
rect 1324 1391 1358 1425
rect 1396 1391 1430 1425
rect 1252 1319 1286 1353
rect 1324 1319 1358 1353
rect 1396 1319 1430 1353
rect 1252 1247 1286 1281
rect 1324 1247 1358 1281
rect 1396 1247 1430 1281
rect 1252 1175 1286 1209
rect 1324 1175 1358 1209
rect 1396 1175 1430 1209
rect 1252 1103 1286 1137
rect 1324 1103 1358 1137
rect 1396 1103 1430 1137
rect 1252 1031 1286 1065
rect 1324 1031 1358 1065
rect 1396 1031 1430 1065
rect 1252 959 1286 993
rect 1324 959 1358 993
rect 1396 959 1430 993
rect 1252 887 1286 921
rect 1324 887 1358 921
rect 1396 887 1430 921
rect 1252 815 1286 849
rect 1324 815 1358 849
rect 1396 815 1430 849
rect 1252 743 1286 777
rect 1324 743 1358 777
rect 1396 743 1430 777
rect 1252 671 1286 705
rect 1324 671 1358 705
rect 1396 671 1430 705
rect 1252 599 1286 633
rect 1324 599 1358 633
rect 1396 599 1430 633
rect 1252 527 1286 561
rect 1324 527 1358 561
rect 1396 527 1430 561
rect 1252 455 1286 489
rect 1324 455 1358 489
rect 1396 455 1430 489
rect 1252 383 1286 417
rect 1324 383 1358 417
rect 1396 383 1430 417
rect 1252 311 1286 345
rect 1324 311 1358 345
rect 1396 311 1430 345
rect 1252 239 1286 273
rect 1324 239 1358 273
rect 1396 239 1430 273
rect 1252 167 1286 201
rect 1324 167 1358 201
rect 1396 167 1430 201
rect 1252 95 1286 129
rect 1324 95 1358 129
rect 1396 95 1430 129
rect 1252 23 1286 57
rect 1324 23 1358 57
rect 1396 23 1430 57
<< poly >>
rect 204 8090 1004 8106
rect 204 8056 227 8090
rect 261 8056 299 8090
rect 333 8056 371 8090
rect 405 8056 443 8090
rect 477 8056 515 8090
rect 549 8056 587 8090
rect 621 8056 659 8090
rect 693 8056 731 8090
rect 765 8056 803 8090
rect 837 8056 875 8090
rect 909 8056 947 8090
rect 981 8056 1004 8090
rect 204 8000 1004 8056
rect 204 -40 1004 0
<< polycont >>
rect 227 8056 261 8090
rect 299 8056 333 8090
rect 371 8056 405 8090
rect 443 8056 477 8090
rect 515 8056 549 8090
rect 587 8056 621 8090
rect 659 8056 693 8090
rect 731 8056 765 8090
rect 803 8056 837 8090
rect 875 8056 909 8090
rect 947 8056 981 8090
<< locali >>
rect 211 8056 227 8090
rect 261 8056 299 8090
rect 333 8056 371 8090
rect 405 8056 443 8090
rect 477 8056 515 8090
rect 549 8056 587 8090
rect 621 8056 659 8090
rect 693 8056 731 8090
rect 765 8056 803 8090
rect 837 8056 875 8090
rect 909 8056 947 8090
rect 981 8056 997 8090
rect 13 7977 191 7993
rect 13 7 191 23
rect 1017 7977 1195 7993
rect 1017 7 1195 23
rect 1252 7977 1430 7993
rect 1286 7943 1324 7977
rect 1358 7943 1396 7977
rect 1252 7905 1430 7943
rect 1286 7871 1324 7905
rect 1358 7871 1396 7905
rect 1252 7833 1430 7871
rect 1286 7799 1324 7833
rect 1358 7799 1396 7833
rect 1252 7761 1430 7799
rect 1286 7727 1324 7761
rect 1358 7727 1396 7761
rect 1252 7689 1430 7727
rect 1286 7655 1324 7689
rect 1358 7655 1396 7689
rect 1252 7617 1430 7655
rect 1286 7583 1324 7617
rect 1358 7583 1396 7617
rect 1252 7545 1430 7583
rect 1286 7511 1324 7545
rect 1358 7511 1396 7545
rect 1252 7473 1430 7511
rect 1286 7439 1324 7473
rect 1358 7439 1396 7473
rect 1252 7401 1430 7439
rect 1286 7367 1324 7401
rect 1358 7367 1396 7401
rect 1252 7329 1430 7367
rect 1286 7295 1324 7329
rect 1358 7295 1396 7329
rect 1252 7257 1430 7295
rect 1286 7223 1324 7257
rect 1358 7223 1396 7257
rect 1252 7185 1430 7223
rect 1286 7151 1324 7185
rect 1358 7151 1396 7185
rect 1252 7113 1430 7151
rect 1286 7079 1324 7113
rect 1358 7079 1396 7113
rect 1252 7041 1430 7079
rect 1286 7007 1324 7041
rect 1358 7007 1396 7041
rect 1252 6969 1430 7007
rect 1286 6935 1324 6969
rect 1358 6935 1396 6969
rect 1252 6897 1430 6935
rect 1286 6863 1324 6897
rect 1358 6863 1396 6897
rect 1252 6825 1430 6863
rect 1286 6791 1324 6825
rect 1358 6791 1396 6825
rect 1252 6753 1430 6791
rect 1286 6719 1324 6753
rect 1358 6719 1396 6753
rect 1252 6681 1430 6719
rect 1286 6647 1324 6681
rect 1358 6647 1396 6681
rect 1252 6609 1430 6647
rect 1286 6575 1324 6609
rect 1358 6575 1396 6609
rect 1252 6537 1430 6575
rect 1286 6503 1324 6537
rect 1358 6503 1396 6537
rect 1252 6465 1430 6503
rect 1286 6431 1324 6465
rect 1358 6431 1396 6465
rect 1252 6393 1430 6431
rect 1286 6359 1324 6393
rect 1358 6359 1396 6393
rect 1252 6321 1430 6359
rect 1286 6287 1324 6321
rect 1358 6287 1396 6321
rect 1252 6249 1430 6287
rect 1286 6215 1324 6249
rect 1358 6215 1396 6249
rect 1252 6177 1430 6215
rect 1286 6143 1324 6177
rect 1358 6143 1396 6177
rect 1252 6105 1430 6143
rect 1286 6071 1324 6105
rect 1358 6071 1396 6105
rect 1252 6033 1430 6071
rect 1286 5999 1324 6033
rect 1358 5999 1396 6033
rect 1252 5961 1430 5999
rect 1286 5927 1324 5961
rect 1358 5927 1396 5961
rect 1252 5889 1430 5927
rect 1286 5855 1324 5889
rect 1358 5855 1396 5889
rect 1252 5817 1430 5855
rect 1286 5783 1324 5817
rect 1358 5783 1396 5817
rect 1252 5745 1430 5783
rect 1286 5711 1324 5745
rect 1358 5711 1396 5745
rect 1252 5673 1430 5711
rect 1286 5639 1324 5673
rect 1358 5639 1396 5673
rect 1252 5601 1430 5639
rect 1286 5567 1324 5601
rect 1358 5567 1396 5601
rect 1252 5529 1430 5567
rect 1286 5495 1324 5529
rect 1358 5495 1396 5529
rect 1252 5457 1430 5495
rect 1286 5423 1324 5457
rect 1358 5423 1396 5457
rect 1252 5385 1430 5423
rect 1286 5351 1324 5385
rect 1358 5351 1396 5385
rect 1252 5313 1430 5351
rect 1286 5279 1324 5313
rect 1358 5279 1396 5313
rect 1252 5241 1430 5279
rect 1286 5207 1324 5241
rect 1358 5207 1396 5241
rect 1252 5169 1430 5207
rect 1286 5135 1324 5169
rect 1358 5135 1396 5169
rect 1252 5097 1430 5135
rect 1286 5063 1324 5097
rect 1358 5063 1396 5097
rect 1252 5025 1430 5063
rect 1286 4991 1324 5025
rect 1358 4991 1396 5025
rect 1252 4953 1430 4991
rect 1286 4919 1324 4953
rect 1358 4919 1396 4953
rect 1252 4881 1430 4919
rect 1286 4847 1324 4881
rect 1358 4847 1396 4881
rect 1252 4809 1430 4847
rect 1286 4775 1324 4809
rect 1358 4775 1396 4809
rect 1252 4737 1430 4775
rect 1286 4703 1324 4737
rect 1358 4703 1396 4737
rect 1252 4665 1430 4703
rect 1286 4631 1324 4665
rect 1358 4631 1396 4665
rect 1252 4593 1430 4631
rect 1286 4559 1324 4593
rect 1358 4559 1396 4593
rect 1252 4521 1430 4559
rect 1286 4487 1324 4521
rect 1358 4487 1396 4521
rect 1252 4449 1430 4487
rect 1286 4415 1324 4449
rect 1358 4415 1396 4449
rect 1252 4377 1430 4415
rect 1286 4343 1324 4377
rect 1358 4343 1396 4377
rect 1252 4305 1430 4343
rect 1286 4271 1324 4305
rect 1358 4271 1396 4305
rect 1252 4233 1430 4271
rect 1286 4199 1324 4233
rect 1358 4199 1396 4233
rect 1252 4161 1430 4199
rect 1286 4127 1324 4161
rect 1358 4127 1396 4161
rect 1252 4089 1430 4127
rect 1286 4055 1324 4089
rect 1358 4055 1396 4089
rect 1252 4017 1430 4055
rect 1286 3983 1324 4017
rect 1358 3983 1396 4017
rect 1252 3945 1430 3983
rect 1286 3911 1324 3945
rect 1358 3911 1396 3945
rect 1252 3873 1430 3911
rect 1286 3839 1324 3873
rect 1358 3839 1396 3873
rect 1252 3801 1430 3839
rect 1286 3767 1324 3801
rect 1358 3767 1396 3801
rect 1252 3729 1430 3767
rect 1286 3695 1324 3729
rect 1358 3695 1396 3729
rect 1252 3657 1430 3695
rect 1286 3623 1324 3657
rect 1358 3623 1396 3657
rect 1252 3585 1430 3623
rect 1286 3551 1324 3585
rect 1358 3551 1396 3585
rect 1252 3513 1430 3551
rect 1286 3479 1324 3513
rect 1358 3479 1396 3513
rect 1252 3441 1430 3479
rect 1286 3407 1324 3441
rect 1358 3407 1396 3441
rect 1252 3369 1430 3407
rect 1286 3335 1324 3369
rect 1358 3335 1396 3369
rect 1252 3297 1430 3335
rect 1286 3263 1324 3297
rect 1358 3263 1396 3297
rect 1252 3225 1430 3263
rect 1286 3191 1324 3225
rect 1358 3191 1396 3225
rect 1252 3153 1430 3191
rect 1286 3119 1324 3153
rect 1358 3119 1396 3153
rect 1252 3081 1430 3119
rect 1286 3047 1324 3081
rect 1358 3047 1396 3081
rect 1252 3009 1430 3047
rect 1286 2975 1324 3009
rect 1358 2975 1396 3009
rect 1252 2937 1430 2975
rect 1286 2903 1324 2937
rect 1358 2903 1396 2937
rect 1252 2865 1430 2903
rect 1286 2831 1324 2865
rect 1358 2831 1396 2865
rect 1252 2793 1430 2831
rect 1286 2759 1324 2793
rect 1358 2759 1396 2793
rect 1252 2721 1430 2759
rect 1286 2687 1324 2721
rect 1358 2687 1396 2721
rect 1252 2649 1430 2687
rect 1286 2615 1324 2649
rect 1358 2615 1396 2649
rect 1252 2577 1430 2615
rect 1286 2543 1324 2577
rect 1358 2543 1396 2577
rect 1252 2505 1430 2543
rect 1286 2471 1324 2505
rect 1358 2471 1396 2505
rect 1252 2433 1430 2471
rect 1286 2399 1324 2433
rect 1358 2399 1396 2433
rect 1252 2361 1430 2399
rect 1286 2327 1324 2361
rect 1358 2327 1396 2361
rect 1252 2289 1430 2327
rect 1286 2255 1324 2289
rect 1358 2255 1396 2289
rect 1252 2217 1430 2255
rect 1286 2183 1324 2217
rect 1358 2183 1396 2217
rect 1252 2145 1430 2183
rect 1286 2111 1324 2145
rect 1358 2111 1396 2145
rect 1252 2073 1430 2111
rect 1286 2039 1324 2073
rect 1358 2039 1396 2073
rect 1252 2001 1430 2039
rect 1286 1967 1324 2001
rect 1358 1967 1396 2001
rect 1252 1929 1430 1967
rect 1286 1895 1324 1929
rect 1358 1895 1396 1929
rect 1252 1857 1430 1895
rect 1286 1823 1324 1857
rect 1358 1823 1396 1857
rect 1252 1785 1430 1823
rect 1286 1751 1324 1785
rect 1358 1751 1396 1785
rect 1252 1713 1430 1751
rect 1286 1679 1324 1713
rect 1358 1679 1396 1713
rect 1252 1641 1430 1679
rect 1286 1607 1324 1641
rect 1358 1607 1396 1641
rect 1252 1569 1430 1607
rect 1286 1535 1324 1569
rect 1358 1535 1396 1569
rect 1252 1497 1430 1535
rect 1286 1463 1324 1497
rect 1358 1463 1396 1497
rect 1252 1425 1430 1463
rect 1286 1391 1324 1425
rect 1358 1391 1396 1425
rect 1252 1353 1430 1391
rect 1286 1319 1324 1353
rect 1358 1319 1396 1353
rect 1252 1281 1430 1319
rect 1286 1247 1324 1281
rect 1358 1247 1396 1281
rect 1252 1209 1430 1247
rect 1286 1175 1324 1209
rect 1358 1175 1396 1209
rect 1252 1137 1430 1175
rect 1286 1103 1324 1137
rect 1358 1103 1396 1137
rect 1252 1065 1430 1103
rect 1286 1031 1324 1065
rect 1358 1031 1396 1065
rect 1252 993 1430 1031
rect 1286 959 1324 993
rect 1358 959 1396 993
rect 1252 921 1430 959
rect 1286 887 1324 921
rect 1358 887 1396 921
rect 1252 849 1430 887
rect 1286 815 1324 849
rect 1358 815 1396 849
rect 1252 777 1430 815
rect 1286 743 1324 777
rect 1358 743 1396 777
rect 1252 705 1430 743
rect 1286 671 1324 705
rect 1358 671 1396 705
rect 1252 633 1430 671
rect 1286 599 1324 633
rect 1358 599 1396 633
rect 1252 561 1430 599
rect 1286 527 1324 561
rect 1358 527 1396 561
rect 1252 489 1430 527
rect 1286 455 1324 489
rect 1358 455 1396 489
rect 1252 417 1430 455
rect 1286 383 1324 417
rect 1358 383 1396 417
rect 1252 345 1430 383
rect 1286 311 1324 345
rect 1358 311 1396 345
rect 1252 273 1430 311
rect 1286 239 1324 273
rect 1358 239 1396 273
rect 1252 201 1430 239
rect 1286 167 1324 201
rect 1358 167 1396 201
rect 1252 129 1430 167
rect 1286 95 1324 129
rect 1358 95 1396 129
rect 1252 57 1430 95
rect 1286 23 1324 57
rect 1358 23 1396 57
rect 1252 7 1430 23
<< viali >>
rect 227 8056 261 8090
rect 299 8056 333 8090
rect 371 8056 405 8090
rect 443 8056 477 8090
rect 515 8056 549 8090
rect 587 8056 621 8090
rect 659 8056 693 8090
rect 731 8056 765 8090
rect 803 8056 837 8090
rect 875 8056 909 8090
rect 947 8056 981 8090
rect 13 7943 47 7977
rect 47 7943 85 7977
rect 85 7943 119 7977
rect 119 7943 157 7977
rect 157 7943 191 7977
rect 13 7905 191 7943
rect 13 7871 47 7905
rect 47 7871 85 7905
rect 85 7871 119 7905
rect 119 7871 157 7905
rect 157 7871 191 7905
rect 13 7833 191 7871
rect 13 7799 47 7833
rect 47 7799 85 7833
rect 85 7799 119 7833
rect 119 7799 157 7833
rect 157 7799 191 7833
rect 13 7761 191 7799
rect 13 7727 47 7761
rect 47 7727 85 7761
rect 85 7727 119 7761
rect 119 7727 157 7761
rect 157 7727 191 7761
rect 13 7689 191 7727
rect 13 7655 47 7689
rect 47 7655 85 7689
rect 85 7655 119 7689
rect 119 7655 157 7689
rect 157 7655 191 7689
rect 13 7617 191 7655
rect 13 7583 47 7617
rect 47 7583 85 7617
rect 85 7583 119 7617
rect 119 7583 157 7617
rect 157 7583 191 7617
rect 13 7545 191 7583
rect 13 7511 47 7545
rect 47 7511 85 7545
rect 85 7511 119 7545
rect 119 7511 157 7545
rect 157 7511 191 7545
rect 13 7473 191 7511
rect 13 7439 47 7473
rect 47 7439 85 7473
rect 85 7439 119 7473
rect 119 7439 157 7473
rect 157 7439 191 7473
rect 13 7401 191 7439
rect 13 7367 47 7401
rect 47 7367 85 7401
rect 85 7367 119 7401
rect 119 7367 157 7401
rect 157 7367 191 7401
rect 13 7329 191 7367
rect 13 7295 47 7329
rect 47 7295 85 7329
rect 85 7295 119 7329
rect 119 7295 157 7329
rect 157 7295 191 7329
rect 13 7257 191 7295
rect 13 7223 47 7257
rect 47 7223 85 7257
rect 85 7223 119 7257
rect 119 7223 157 7257
rect 157 7223 191 7257
rect 13 7185 191 7223
rect 13 7151 47 7185
rect 47 7151 85 7185
rect 85 7151 119 7185
rect 119 7151 157 7185
rect 157 7151 191 7185
rect 13 7113 191 7151
rect 13 7079 47 7113
rect 47 7079 85 7113
rect 85 7079 119 7113
rect 119 7079 157 7113
rect 157 7079 191 7113
rect 13 7041 191 7079
rect 13 7007 47 7041
rect 47 7007 85 7041
rect 85 7007 119 7041
rect 119 7007 157 7041
rect 157 7007 191 7041
rect 13 6969 191 7007
rect 13 6935 47 6969
rect 47 6935 85 6969
rect 85 6935 119 6969
rect 119 6935 157 6969
rect 157 6935 191 6969
rect 13 6897 191 6935
rect 13 6863 47 6897
rect 47 6863 85 6897
rect 85 6863 119 6897
rect 119 6863 157 6897
rect 157 6863 191 6897
rect 13 6825 191 6863
rect 13 6791 47 6825
rect 47 6791 85 6825
rect 85 6791 119 6825
rect 119 6791 157 6825
rect 157 6791 191 6825
rect 13 6753 191 6791
rect 13 6719 47 6753
rect 47 6719 85 6753
rect 85 6719 119 6753
rect 119 6719 157 6753
rect 157 6719 191 6753
rect 13 6681 191 6719
rect 13 6647 47 6681
rect 47 6647 85 6681
rect 85 6647 119 6681
rect 119 6647 157 6681
rect 157 6647 191 6681
rect 13 6609 191 6647
rect 13 6575 47 6609
rect 47 6575 85 6609
rect 85 6575 119 6609
rect 119 6575 157 6609
rect 157 6575 191 6609
rect 13 6537 191 6575
rect 13 6503 47 6537
rect 47 6503 85 6537
rect 85 6503 119 6537
rect 119 6503 157 6537
rect 157 6503 191 6537
rect 13 6465 191 6503
rect 13 6431 47 6465
rect 47 6431 85 6465
rect 85 6431 119 6465
rect 119 6431 157 6465
rect 157 6431 191 6465
rect 13 6393 191 6431
rect 13 6359 47 6393
rect 47 6359 85 6393
rect 85 6359 119 6393
rect 119 6359 157 6393
rect 157 6359 191 6393
rect 13 6321 191 6359
rect 13 6287 47 6321
rect 47 6287 85 6321
rect 85 6287 119 6321
rect 119 6287 157 6321
rect 157 6287 191 6321
rect 13 6249 191 6287
rect 13 6215 47 6249
rect 47 6215 85 6249
rect 85 6215 119 6249
rect 119 6215 157 6249
rect 157 6215 191 6249
rect 13 6177 191 6215
rect 13 6143 47 6177
rect 47 6143 85 6177
rect 85 6143 119 6177
rect 119 6143 157 6177
rect 157 6143 191 6177
rect 13 6105 191 6143
rect 13 6071 47 6105
rect 47 6071 85 6105
rect 85 6071 119 6105
rect 119 6071 157 6105
rect 157 6071 191 6105
rect 13 6033 191 6071
rect 13 5999 47 6033
rect 47 5999 85 6033
rect 85 5999 119 6033
rect 119 5999 157 6033
rect 157 5999 191 6033
rect 13 5961 191 5999
rect 13 5927 47 5961
rect 47 5927 85 5961
rect 85 5927 119 5961
rect 119 5927 157 5961
rect 157 5927 191 5961
rect 13 5889 191 5927
rect 13 5855 47 5889
rect 47 5855 85 5889
rect 85 5855 119 5889
rect 119 5855 157 5889
rect 157 5855 191 5889
rect 13 5817 191 5855
rect 13 5783 47 5817
rect 47 5783 85 5817
rect 85 5783 119 5817
rect 119 5783 157 5817
rect 157 5783 191 5817
rect 13 5745 191 5783
rect 13 5711 47 5745
rect 47 5711 85 5745
rect 85 5711 119 5745
rect 119 5711 157 5745
rect 157 5711 191 5745
rect 13 5673 191 5711
rect 13 5639 47 5673
rect 47 5639 85 5673
rect 85 5639 119 5673
rect 119 5639 157 5673
rect 157 5639 191 5673
rect 13 5601 191 5639
rect 13 5567 47 5601
rect 47 5567 85 5601
rect 85 5567 119 5601
rect 119 5567 157 5601
rect 157 5567 191 5601
rect 13 5529 191 5567
rect 13 5495 47 5529
rect 47 5495 85 5529
rect 85 5495 119 5529
rect 119 5495 157 5529
rect 157 5495 191 5529
rect 13 5457 191 5495
rect 13 5423 47 5457
rect 47 5423 85 5457
rect 85 5423 119 5457
rect 119 5423 157 5457
rect 157 5423 191 5457
rect 13 5385 191 5423
rect 13 5351 47 5385
rect 47 5351 85 5385
rect 85 5351 119 5385
rect 119 5351 157 5385
rect 157 5351 191 5385
rect 13 5313 191 5351
rect 13 5279 47 5313
rect 47 5279 85 5313
rect 85 5279 119 5313
rect 119 5279 157 5313
rect 157 5279 191 5313
rect 13 5241 191 5279
rect 13 5207 47 5241
rect 47 5207 85 5241
rect 85 5207 119 5241
rect 119 5207 157 5241
rect 157 5207 191 5241
rect 13 5169 191 5207
rect 13 5135 47 5169
rect 47 5135 85 5169
rect 85 5135 119 5169
rect 119 5135 157 5169
rect 157 5135 191 5169
rect 13 5097 191 5135
rect 13 5063 47 5097
rect 47 5063 85 5097
rect 85 5063 119 5097
rect 119 5063 157 5097
rect 157 5063 191 5097
rect 13 5025 191 5063
rect 13 4991 47 5025
rect 47 4991 85 5025
rect 85 4991 119 5025
rect 119 4991 157 5025
rect 157 4991 191 5025
rect 13 4953 191 4991
rect 13 4919 47 4953
rect 47 4919 85 4953
rect 85 4919 119 4953
rect 119 4919 157 4953
rect 157 4919 191 4953
rect 13 4881 191 4919
rect 13 4847 47 4881
rect 47 4847 85 4881
rect 85 4847 119 4881
rect 119 4847 157 4881
rect 157 4847 191 4881
rect 13 4809 191 4847
rect 13 4775 47 4809
rect 47 4775 85 4809
rect 85 4775 119 4809
rect 119 4775 157 4809
rect 157 4775 191 4809
rect 13 4737 191 4775
rect 13 4703 47 4737
rect 47 4703 85 4737
rect 85 4703 119 4737
rect 119 4703 157 4737
rect 157 4703 191 4737
rect 13 4665 191 4703
rect 13 4631 47 4665
rect 47 4631 85 4665
rect 85 4631 119 4665
rect 119 4631 157 4665
rect 157 4631 191 4665
rect 13 4593 191 4631
rect 13 4559 47 4593
rect 47 4559 85 4593
rect 85 4559 119 4593
rect 119 4559 157 4593
rect 157 4559 191 4593
rect 13 4521 191 4559
rect 13 4487 47 4521
rect 47 4487 85 4521
rect 85 4487 119 4521
rect 119 4487 157 4521
rect 157 4487 191 4521
rect 13 4449 191 4487
rect 13 4415 47 4449
rect 47 4415 85 4449
rect 85 4415 119 4449
rect 119 4415 157 4449
rect 157 4415 191 4449
rect 13 4377 191 4415
rect 13 4343 47 4377
rect 47 4343 85 4377
rect 85 4343 119 4377
rect 119 4343 157 4377
rect 157 4343 191 4377
rect 13 4305 191 4343
rect 13 4271 47 4305
rect 47 4271 85 4305
rect 85 4271 119 4305
rect 119 4271 157 4305
rect 157 4271 191 4305
rect 13 4233 191 4271
rect 13 4199 47 4233
rect 47 4199 85 4233
rect 85 4199 119 4233
rect 119 4199 157 4233
rect 157 4199 191 4233
rect 13 4161 191 4199
rect 13 4127 47 4161
rect 47 4127 85 4161
rect 85 4127 119 4161
rect 119 4127 157 4161
rect 157 4127 191 4161
rect 13 4089 191 4127
rect 13 4055 47 4089
rect 47 4055 85 4089
rect 85 4055 119 4089
rect 119 4055 157 4089
rect 157 4055 191 4089
rect 13 4017 191 4055
rect 13 3983 47 4017
rect 47 3983 85 4017
rect 85 3983 119 4017
rect 119 3983 157 4017
rect 157 3983 191 4017
rect 13 3945 191 3983
rect 13 3911 47 3945
rect 47 3911 85 3945
rect 85 3911 119 3945
rect 119 3911 157 3945
rect 157 3911 191 3945
rect 13 3873 191 3911
rect 13 3839 47 3873
rect 47 3839 85 3873
rect 85 3839 119 3873
rect 119 3839 157 3873
rect 157 3839 191 3873
rect 13 3801 191 3839
rect 13 3767 47 3801
rect 47 3767 85 3801
rect 85 3767 119 3801
rect 119 3767 157 3801
rect 157 3767 191 3801
rect 13 3729 191 3767
rect 13 3695 47 3729
rect 47 3695 85 3729
rect 85 3695 119 3729
rect 119 3695 157 3729
rect 157 3695 191 3729
rect 13 3657 191 3695
rect 13 3623 47 3657
rect 47 3623 85 3657
rect 85 3623 119 3657
rect 119 3623 157 3657
rect 157 3623 191 3657
rect 13 3585 191 3623
rect 13 3551 47 3585
rect 47 3551 85 3585
rect 85 3551 119 3585
rect 119 3551 157 3585
rect 157 3551 191 3585
rect 13 3513 191 3551
rect 13 3479 47 3513
rect 47 3479 85 3513
rect 85 3479 119 3513
rect 119 3479 157 3513
rect 157 3479 191 3513
rect 13 3441 191 3479
rect 13 3407 47 3441
rect 47 3407 85 3441
rect 85 3407 119 3441
rect 119 3407 157 3441
rect 157 3407 191 3441
rect 13 3369 191 3407
rect 13 3335 47 3369
rect 47 3335 85 3369
rect 85 3335 119 3369
rect 119 3335 157 3369
rect 157 3335 191 3369
rect 13 3297 191 3335
rect 13 3263 47 3297
rect 47 3263 85 3297
rect 85 3263 119 3297
rect 119 3263 157 3297
rect 157 3263 191 3297
rect 13 3225 191 3263
rect 13 3191 47 3225
rect 47 3191 85 3225
rect 85 3191 119 3225
rect 119 3191 157 3225
rect 157 3191 191 3225
rect 13 3153 191 3191
rect 13 3119 47 3153
rect 47 3119 85 3153
rect 85 3119 119 3153
rect 119 3119 157 3153
rect 157 3119 191 3153
rect 13 3081 191 3119
rect 13 3047 47 3081
rect 47 3047 85 3081
rect 85 3047 119 3081
rect 119 3047 157 3081
rect 157 3047 191 3081
rect 13 3009 191 3047
rect 13 2975 47 3009
rect 47 2975 85 3009
rect 85 2975 119 3009
rect 119 2975 157 3009
rect 157 2975 191 3009
rect 13 2937 191 2975
rect 13 2903 47 2937
rect 47 2903 85 2937
rect 85 2903 119 2937
rect 119 2903 157 2937
rect 157 2903 191 2937
rect 13 2865 191 2903
rect 13 2831 47 2865
rect 47 2831 85 2865
rect 85 2831 119 2865
rect 119 2831 157 2865
rect 157 2831 191 2865
rect 13 2793 191 2831
rect 13 2759 47 2793
rect 47 2759 85 2793
rect 85 2759 119 2793
rect 119 2759 157 2793
rect 157 2759 191 2793
rect 13 2721 191 2759
rect 13 2687 47 2721
rect 47 2687 85 2721
rect 85 2687 119 2721
rect 119 2687 157 2721
rect 157 2687 191 2721
rect 13 2649 191 2687
rect 13 2615 47 2649
rect 47 2615 85 2649
rect 85 2615 119 2649
rect 119 2615 157 2649
rect 157 2615 191 2649
rect 13 2577 191 2615
rect 13 2543 47 2577
rect 47 2543 85 2577
rect 85 2543 119 2577
rect 119 2543 157 2577
rect 157 2543 191 2577
rect 13 2505 191 2543
rect 13 2471 47 2505
rect 47 2471 85 2505
rect 85 2471 119 2505
rect 119 2471 157 2505
rect 157 2471 191 2505
rect 13 2433 191 2471
rect 13 2399 47 2433
rect 47 2399 85 2433
rect 85 2399 119 2433
rect 119 2399 157 2433
rect 157 2399 191 2433
rect 13 2361 191 2399
rect 13 2327 47 2361
rect 47 2327 85 2361
rect 85 2327 119 2361
rect 119 2327 157 2361
rect 157 2327 191 2361
rect 13 2289 191 2327
rect 13 2255 47 2289
rect 47 2255 85 2289
rect 85 2255 119 2289
rect 119 2255 157 2289
rect 157 2255 191 2289
rect 13 2217 191 2255
rect 13 2183 47 2217
rect 47 2183 85 2217
rect 85 2183 119 2217
rect 119 2183 157 2217
rect 157 2183 191 2217
rect 13 2145 191 2183
rect 13 2111 47 2145
rect 47 2111 85 2145
rect 85 2111 119 2145
rect 119 2111 157 2145
rect 157 2111 191 2145
rect 13 2073 191 2111
rect 13 2039 47 2073
rect 47 2039 85 2073
rect 85 2039 119 2073
rect 119 2039 157 2073
rect 157 2039 191 2073
rect 13 2001 191 2039
rect 13 1967 47 2001
rect 47 1967 85 2001
rect 85 1967 119 2001
rect 119 1967 157 2001
rect 157 1967 191 2001
rect 13 1929 191 1967
rect 13 1895 47 1929
rect 47 1895 85 1929
rect 85 1895 119 1929
rect 119 1895 157 1929
rect 157 1895 191 1929
rect 13 1857 191 1895
rect 13 1823 47 1857
rect 47 1823 85 1857
rect 85 1823 119 1857
rect 119 1823 157 1857
rect 157 1823 191 1857
rect 13 1785 191 1823
rect 13 1751 47 1785
rect 47 1751 85 1785
rect 85 1751 119 1785
rect 119 1751 157 1785
rect 157 1751 191 1785
rect 13 1713 191 1751
rect 13 1679 47 1713
rect 47 1679 85 1713
rect 85 1679 119 1713
rect 119 1679 157 1713
rect 157 1679 191 1713
rect 13 1641 191 1679
rect 13 1607 47 1641
rect 47 1607 85 1641
rect 85 1607 119 1641
rect 119 1607 157 1641
rect 157 1607 191 1641
rect 13 1569 191 1607
rect 13 1535 47 1569
rect 47 1535 85 1569
rect 85 1535 119 1569
rect 119 1535 157 1569
rect 157 1535 191 1569
rect 13 1497 191 1535
rect 13 1463 47 1497
rect 47 1463 85 1497
rect 85 1463 119 1497
rect 119 1463 157 1497
rect 157 1463 191 1497
rect 13 1425 191 1463
rect 13 1391 47 1425
rect 47 1391 85 1425
rect 85 1391 119 1425
rect 119 1391 157 1425
rect 157 1391 191 1425
rect 13 1353 191 1391
rect 13 1319 47 1353
rect 47 1319 85 1353
rect 85 1319 119 1353
rect 119 1319 157 1353
rect 157 1319 191 1353
rect 13 1281 191 1319
rect 13 1247 47 1281
rect 47 1247 85 1281
rect 85 1247 119 1281
rect 119 1247 157 1281
rect 157 1247 191 1281
rect 13 1209 191 1247
rect 13 1175 47 1209
rect 47 1175 85 1209
rect 85 1175 119 1209
rect 119 1175 157 1209
rect 157 1175 191 1209
rect 13 1137 191 1175
rect 13 1103 47 1137
rect 47 1103 85 1137
rect 85 1103 119 1137
rect 119 1103 157 1137
rect 157 1103 191 1137
rect 13 1065 191 1103
rect 13 1031 47 1065
rect 47 1031 85 1065
rect 85 1031 119 1065
rect 119 1031 157 1065
rect 157 1031 191 1065
rect 13 993 191 1031
rect 13 959 47 993
rect 47 959 85 993
rect 85 959 119 993
rect 119 959 157 993
rect 157 959 191 993
rect 13 921 191 959
rect 13 887 47 921
rect 47 887 85 921
rect 85 887 119 921
rect 119 887 157 921
rect 157 887 191 921
rect 13 849 191 887
rect 13 815 47 849
rect 47 815 85 849
rect 85 815 119 849
rect 119 815 157 849
rect 157 815 191 849
rect 13 777 191 815
rect 13 743 47 777
rect 47 743 85 777
rect 85 743 119 777
rect 119 743 157 777
rect 157 743 191 777
rect 13 705 191 743
rect 13 671 47 705
rect 47 671 85 705
rect 85 671 119 705
rect 119 671 157 705
rect 157 671 191 705
rect 13 633 191 671
rect 13 599 47 633
rect 47 599 85 633
rect 85 599 119 633
rect 119 599 157 633
rect 157 599 191 633
rect 13 561 191 599
rect 13 527 47 561
rect 47 527 85 561
rect 85 527 119 561
rect 119 527 157 561
rect 157 527 191 561
rect 13 489 191 527
rect 13 455 47 489
rect 47 455 85 489
rect 85 455 119 489
rect 119 455 157 489
rect 157 455 191 489
rect 13 417 191 455
rect 13 383 47 417
rect 47 383 85 417
rect 85 383 119 417
rect 119 383 157 417
rect 157 383 191 417
rect 13 345 191 383
rect 13 311 47 345
rect 47 311 85 345
rect 85 311 119 345
rect 119 311 157 345
rect 157 311 191 345
rect 13 273 191 311
rect 13 239 47 273
rect 47 239 85 273
rect 85 239 119 273
rect 119 239 157 273
rect 157 239 191 273
rect 13 201 191 239
rect 13 167 47 201
rect 47 167 85 201
rect 85 167 119 201
rect 119 167 157 201
rect 157 167 191 201
rect 13 129 191 167
rect 13 95 47 129
rect 47 95 85 129
rect 85 95 119 129
rect 119 95 157 129
rect 157 95 191 129
rect 13 57 191 95
rect 13 23 47 57
rect 47 23 85 57
rect 85 23 119 57
rect 119 23 157 57
rect 157 23 191 57
rect 1017 7943 1051 7977
rect 1051 7943 1089 7977
rect 1089 7943 1123 7977
rect 1123 7943 1161 7977
rect 1161 7943 1195 7977
rect 1017 7905 1195 7943
rect 1017 7871 1051 7905
rect 1051 7871 1089 7905
rect 1089 7871 1123 7905
rect 1123 7871 1161 7905
rect 1161 7871 1195 7905
rect 1017 7833 1195 7871
rect 1017 7799 1051 7833
rect 1051 7799 1089 7833
rect 1089 7799 1123 7833
rect 1123 7799 1161 7833
rect 1161 7799 1195 7833
rect 1017 7761 1195 7799
rect 1017 7727 1051 7761
rect 1051 7727 1089 7761
rect 1089 7727 1123 7761
rect 1123 7727 1161 7761
rect 1161 7727 1195 7761
rect 1017 7689 1195 7727
rect 1017 7655 1051 7689
rect 1051 7655 1089 7689
rect 1089 7655 1123 7689
rect 1123 7655 1161 7689
rect 1161 7655 1195 7689
rect 1017 7617 1195 7655
rect 1017 7583 1051 7617
rect 1051 7583 1089 7617
rect 1089 7583 1123 7617
rect 1123 7583 1161 7617
rect 1161 7583 1195 7617
rect 1017 7545 1195 7583
rect 1017 7511 1051 7545
rect 1051 7511 1089 7545
rect 1089 7511 1123 7545
rect 1123 7511 1161 7545
rect 1161 7511 1195 7545
rect 1017 7473 1195 7511
rect 1017 7439 1051 7473
rect 1051 7439 1089 7473
rect 1089 7439 1123 7473
rect 1123 7439 1161 7473
rect 1161 7439 1195 7473
rect 1017 7401 1195 7439
rect 1017 7367 1051 7401
rect 1051 7367 1089 7401
rect 1089 7367 1123 7401
rect 1123 7367 1161 7401
rect 1161 7367 1195 7401
rect 1017 7329 1195 7367
rect 1017 7295 1051 7329
rect 1051 7295 1089 7329
rect 1089 7295 1123 7329
rect 1123 7295 1161 7329
rect 1161 7295 1195 7329
rect 1017 7257 1195 7295
rect 1017 7223 1051 7257
rect 1051 7223 1089 7257
rect 1089 7223 1123 7257
rect 1123 7223 1161 7257
rect 1161 7223 1195 7257
rect 1017 7185 1195 7223
rect 1017 7151 1051 7185
rect 1051 7151 1089 7185
rect 1089 7151 1123 7185
rect 1123 7151 1161 7185
rect 1161 7151 1195 7185
rect 1017 7113 1195 7151
rect 1017 7079 1051 7113
rect 1051 7079 1089 7113
rect 1089 7079 1123 7113
rect 1123 7079 1161 7113
rect 1161 7079 1195 7113
rect 1017 7041 1195 7079
rect 1017 7007 1051 7041
rect 1051 7007 1089 7041
rect 1089 7007 1123 7041
rect 1123 7007 1161 7041
rect 1161 7007 1195 7041
rect 1017 6969 1195 7007
rect 1017 6935 1051 6969
rect 1051 6935 1089 6969
rect 1089 6935 1123 6969
rect 1123 6935 1161 6969
rect 1161 6935 1195 6969
rect 1017 6897 1195 6935
rect 1017 6863 1051 6897
rect 1051 6863 1089 6897
rect 1089 6863 1123 6897
rect 1123 6863 1161 6897
rect 1161 6863 1195 6897
rect 1017 6825 1195 6863
rect 1017 6791 1051 6825
rect 1051 6791 1089 6825
rect 1089 6791 1123 6825
rect 1123 6791 1161 6825
rect 1161 6791 1195 6825
rect 1017 6753 1195 6791
rect 1017 6719 1051 6753
rect 1051 6719 1089 6753
rect 1089 6719 1123 6753
rect 1123 6719 1161 6753
rect 1161 6719 1195 6753
rect 1017 6681 1195 6719
rect 1017 6647 1051 6681
rect 1051 6647 1089 6681
rect 1089 6647 1123 6681
rect 1123 6647 1161 6681
rect 1161 6647 1195 6681
rect 1017 6609 1195 6647
rect 1017 6575 1051 6609
rect 1051 6575 1089 6609
rect 1089 6575 1123 6609
rect 1123 6575 1161 6609
rect 1161 6575 1195 6609
rect 1017 6537 1195 6575
rect 1017 6503 1051 6537
rect 1051 6503 1089 6537
rect 1089 6503 1123 6537
rect 1123 6503 1161 6537
rect 1161 6503 1195 6537
rect 1017 6465 1195 6503
rect 1017 6431 1051 6465
rect 1051 6431 1089 6465
rect 1089 6431 1123 6465
rect 1123 6431 1161 6465
rect 1161 6431 1195 6465
rect 1017 6393 1195 6431
rect 1017 6359 1051 6393
rect 1051 6359 1089 6393
rect 1089 6359 1123 6393
rect 1123 6359 1161 6393
rect 1161 6359 1195 6393
rect 1017 6321 1195 6359
rect 1017 6287 1051 6321
rect 1051 6287 1089 6321
rect 1089 6287 1123 6321
rect 1123 6287 1161 6321
rect 1161 6287 1195 6321
rect 1017 6249 1195 6287
rect 1017 6215 1051 6249
rect 1051 6215 1089 6249
rect 1089 6215 1123 6249
rect 1123 6215 1161 6249
rect 1161 6215 1195 6249
rect 1017 6177 1195 6215
rect 1017 6143 1051 6177
rect 1051 6143 1089 6177
rect 1089 6143 1123 6177
rect 1123 6143 1161 6177
rect 1161 6143 1195 6177
rect 1017 6105 1195 6143
rect 1017 6071 1051 6105
rect 1051 6071 1089 6105
rect 1089 6071 1123 6105
rect 1123 6071 1161 6105
rect 1161 6071 1195 6105
rect 1017 6033 1195 6071
rect 1017 5999 1051 6033
rect 1051 5999 1089 6033
rect 1089 5999 1123 6033
rect 1123 5999 1161 6033
rect 1161 5999 1195 6033
rect 1017 5961 1195 5999
rect 1017 5927 1051 5961
rect 1051 5927 1089 5961
rect 1089 5927 1123 5961
rect 1123 5927 1161 5961
rect 1161 5927 1195 5961
rect 1017 5889 1195 5927
rect 1017 5855 1051 5889
rect 1051 5855 1089 5889
rect 1089 5855 1123 5889
rect 1123 5855 1161 5889
rect 1161 5855 1195 5889
rect 1017 5817 1195 5855
rect 1017 5783 1051 5817
rect 1051 5783 1089 5817
rect 1089 5783 1123 5817
rect 1123 5783 1161 5817
rect 1161 5783 1195 5817
rect 1017 5745 1195 5783
rect 1017 5711 1051 5745
rect 1051 5711 1089 5745
rect 1089 5711 1123 5745
rect 1123 5711 1161 5745
rect 1161 5711 1195 5745
rect 1017 5673 1195 5711
rect 1017 5639 1051 5673
rect 1051 5639 1089 5673
rect 1089 5639 1123 5673
rect 1123 5639 1161 5673
rect 1161 5639 1195 5673
rect 1017 5601 1195 5639
rect 1017 5567 1051 5601
rect 1051 5567 1089 5601
rect 1089 5567 1123 5601
rect 1123 5567 1161 5601
rect 1161 5567 1195 5601
rect 1017 5529 1195 5567
rect 1017 5495 1051 5529
rect 1051 5495 1089 5529
rect 1089 5495 1123 5529
rect 1123 5495 1161 5529
rect 1161 5495 1195 5529
rect 1017 5457 1195 5495
rect 1017 5423 1051 5457
rect 1051 5423 1089 5457
rect 1089 5423 1123 5457
rect 1123 5423 1161 5457
rect 1161 5423 1195 5457
rect 1017 5385 1195 5423
rect 1017 5351 1051 5385
rect 1051 5351 1089 5385
rect 1089 5351 1123 5385
rect 1123 5351 1161 5385
rect 1161 5351 1195 5385
rect 1017 5313 1195 5351
rect 1017 5279 1051 5313
rect 1051 5279 1089 5313
rect 1089 5279 1123 5313
rect 1123 5279 1161 5313
rect 1161 5279 1195 5313
rect 1017 5241 1195 5279
rect 1017 5207 1051 5241
rect 1051 5207 1089 5241
rect 1089 5207 1123 5241
rect 1123 5207 1161 5241
rect 1161 5207 1195 5241
rect 1017 5169 1195 5207
rect 1017 5135 1051 5169
rect 1051 5135 1089 5169
rect 1089 5135 1123 5169
rect 1123 5135 1161 5169
rect 1161 5135 1195 5169
rect 1017 5097 1195 5135
rect 1017 5063 1051 5097
rect 1051 5063 1089 5097
rect 1089 5063 1123 5097
rect 1123 5063 1161 5097
rect 1161 5063 1195 5097
rect 1017 5025 1195 5063
rect 1017 4991 1051 5025
rect 1051 4991 1089 5025
rect 1089 4991 1123 5025
rect 1123 4991 1161 5025
rect 1161 4991 1195 5025
rect 1017 4953 1195 4991
rect 1017 4919 1051 4953
rect 1051 4919 1089 4953
rect 1089 4919 1123 4953
rect 1123 4919 1161 4953
rect 1161 4919 1195 4953
rect 1017 4881 1195 4919
rect 1017 4847 1051 4881
rect 1051 4847 1089 4881
rect 1089 4847 1123 4881
rect 1123 4847 1161 4881
rect 1161 4847 1195 4881
rect 1017 4809 1195 4847
rect 1017 4775 1051 4809
rect 1051 4775 1089 4809
rect 1089 4775 1123 4809
rect 1123 4775 1161 4809
rect 1161 4775 1195 4809
rect 1017 4737 1195 4775
rect 1017 4703 1051 4737
rect 1051 4703 1089 4737
rect 1089 4703 1123 4737
rect 1123 4703 1161 4737
rect 1161 4703 1195 4737
rect 1017 4665 1195 4703
rect 1017 4631 1051 4665
rect 1051 4631 1089 4665
rect 1089 4631 1123 4665
rect 1123 4631 1161 4665
rect 1161 4631 1195 4665
rect 1017 4593 1195 4631
rect 1017 4559 1051 4593
rect 1051 4559 1089 4593
rect 1089 4559 1123 4593
rect 1123 4559 1161 4593
rect 1161 4559 1195 4593
rect 1017 4521 1195 4559
rect 1017 4487 1051 4521
rect 1051 4487 1089 4521
rect 1089 4487 1123 4521
rect 1123 4487 1161 4521
rect 1161 4487 1195 4521
rect 1017 4449 1195 4487
rect 1017 4415 1051 4449
rect 1051 4415 1089 4449
rect 1089 4415 1123 4449
rect 1123 4415 1161 4449
rect 1161 4415 1195 4449
rect 1017 4377 1195 4415
rect 1017 4343 1051 4377
rect 1051 4343 1089 4377
rect 1089 4343 1123 4377
rect 1123 4343 1161 4377
rect 1161 4343 1195 4377
rect 1017 4305 1195 4343
rect 1017 4271 1051 4305
rect 1051 4271 1089 4305
rect 1089 4271 1123 4305
rect 1123 4271 1161 4305
rect 1161 4271 1195 4305
rect 1017 4233 1195 4271
rect 1017 4199 1051 4233
rect 1051 4199 1089 4233
rect 1089 4199 1123 4233
rect 1123 4199 1161 4233
rect 1161 4199 1195 4233
rect 1017 4161 1195 4199
rect 1017 4127 1051 4161
rect 1051 4127 1089 4161
rect 1089 4127 1123 4161
rect 1123 4127 1161 4161
rect 1161 4127 1195 4161
rect 1017 4089 1195 4127
rect 1017 4055 1051 4089
rect 1051 4055 1089 4089
rect 1089 4055 1123 4089
rect 1123 4055 1161 4089
rect 1161 4055 1195 4089
rect 1017 4017 1195 4055
rect 1017 3983 1051 4017
rect 1051 3983 1089 4017
rect 1089 3983 1123 4017
rect 1123 3983 1161 4017
rect 1161 3983 1195 4017
rect 1017 3945 1195 3983
rect 1017 3911 1051 3945
rect 1051 3911 1089 3945
rect 1089 3911 1123 3945
rect 1123 3911 1161 3945
rect 1161 3911 1195 3945
rect 1017 3873 1195 3911
rect 1017 3839 1051 3873
rect 1051 3839 1089 3873
rect 1089 3839 1123 3873
rect 1123 3839 1161 3873
rect 1161 3839 1195 3873
rect 1017 3801 1195 3839
rect 1017 3767 1051 3801
rect 1051 3767 1089 3801
rect 1089 3767 1123 3801
rect 1123 3767 1161 3801
rect 1161 3767 1195 3801
rect 1017 3729 1195 3767
rect 1017 3695 1051 3729
rect 1051 3695 1089 3729
rect 1089 3695 1123 3729
rect 1123 3695 1161 3729
rect 1161 3695 1195 3729
rect 1017 3657 1195 3695
rect 1017 3623 1051 3657
rect 1051 3623 1089 3657
rect 1089 3623 1123 3657
rect 1123 3623 1161 3657
rect 1161 3623 1195 3657
rect 1017 3585 1195 3623
rect 1017 3551 1051 3585
rect 1051 3551 1089 3585
rect 1089 3551 1123 3585
rect 1123 3551 1161 3585
rect 1161 3551 1195 3585
rect 1017 3513 1195 3551
rect 1017 3479 1051 3513
rect 1051 3479 1089 3513
rect 1089 3479 1123 3513
rect 1123 3479 1161 3513
rect 1161 3479 1195 3513
rect 1017 3441 1195 3479
rect 1017 3407 1051 3441
rect 1051 3407 1089 3441
rect 1089 3407 1123 3441
rect 1123 3407 1161 3441
rect 1161 3407 1195 3441
rect 1017 3369 1195 3407
rect 1017 3335 1051 3369
rect 1051 3335 1089 3369
rect 1089 3335 1123 3369
rect 1123 3335 1161 3369
rect 1161 3335 1195 3369
rect 1017 3297 1195 3335
rect 1017 3263 1051 3297
rect 1051 3263 1089 3297
rect 1089 3263 1123 3297
rect 1123 3263 1161 3297
rect 1161 3263 1195 3297
rect 1017 3225 1195 3263
rect 1017 3191 1051 3225
rect 1051 3191 1089 3225
rect 1089 3191 1123 3225
rect 1123 3191 1161 3225
rect 1161 3191 1195 3225
rect 1017 3153 1195 3191
rect 1017 3119 1051 3153
rect 1051 3119 1089 3153
rect 1089 3119 1123 3153
rect 1123 3119 1161 3153
rect 1161 3119 1195 3153
rect 1017 3081 1195 3119
rect 1017 3047 1051 3081
rect 1051 3047 1089 3081
rect 1089 3047 1123 3081
rect 1123 3047 1161 3081
rect 1161 3047 1195 3081
rect 1017 3009 1195 3047
rect 1017 2975 1051 3009
rect 1051 2975 1089 3009
rect 1089 2975 1123 3009
rect 1123 2975 1161 3009
rect 1161 2975 1195 3009
rect 1017 2937 1195 2975
rect 1017 2903 1051 2937
rect 1051 2903 1089 2937
rect 1089 2903 1123 2937
rect 1123 2903 1161 2937
rect 1161 2903 1195 2937
rect 1017 2865 1195 2903
rect 1017 2831 1051 2865
rect 1051 2831 1089 2865
rect 1089 2831 1123 2865
rect 1123 2831 1161 2865
rect 1161 2831 1195 2865
rect 1017 2793 1195 2831
rect 1017 2759 1051 2793
rect 1051 2759 1089 2793
rect 1089 2759 1123 2793
rect 1123 2759 1161 2793
rect 1161 2759 1195 2793
rect 1017 2721 1195 2759
rect 1017 2687 1051 2721
rect 1051 2687 1089 2721
rect 1089 2687 1123 2721
rect 1123 2687 1161 2721
rect 1161 2687 1195 2721
rect 1017 2649 1195 2687
rect 1017 2615 1051 2649
rect 1051 2615 1089 2649
rect 1089 2615 1123 2649
rect 1123 2615 1161 2649
rect 1161 2615 1195 2649
rect 1017 2577 1195 2615
rect 1017 2543 1051 2577
rect 1051 2543 1089 2577
rect 1089 2543 1123 2577
rect 1123 2543 1161 2577
rect 1161 2543 1195 2577
rect 1017 2505 1195 2543
rect 1017 2471 1051 2505
rect 1051 2471 1089 2505
rect 1089 2471 1123 2505
rect 1123 2471 1161 2505
rect 1161 2471 1195 2505
rect 1017 2433 1195 2471
rect 1017 2399 1051 2433
rect 1051 2399 1089 2433
rect 1089 2399 1123 2433
rect 1123 2399 1161 2433
rect 1161 2399 1195 2433
rect 1017 2361 1195 2399
rect 1017 2327 1051 2361
rect 1051 2327 1089 2361
rect 1089 2327 1123 2361
rect 1123 2327 1161 2361
rect 1161 2327 1195 2361
rect 1017 2289 1195 2327
rect 1017 2255 1051 2289
rect 1051 2255 1089 2289
rect 1089 2255 1123 2289
rect 1123 2255 1161 2289
rect 1161 2255 1195 2289
rect 1017 2217 1195 2255
rect 1017 2183 1051 2217
rect 1051 2183 1089 2217
rect 1089 2183 1123 2217
rect 1123 2183 1161 2217
rect 1161 2183 1195 2217
rect 1017 2145 1195 2183
rect 1017 2111 1051 2145
rect 1051 2111 1089 2145
rect 1089 2111 1123 2145
rect 1123 2111 1161 2145
rect 1161 2111 1195 2145
rect 1017 2073 1195 2111
rect 1017 2039 1051 2073
rect 1051 2039 1089 2073
rect 1089 2039 1123 2073
rect 1123 2039 1161 2073
rect 1161 2039 1195 2073
rect 1017 2001 1195 2039
rect 1017 1967 1051 2001
rect 1051 1967 1089 2001
rect 1089 1967 1123 2001
rect 1123 1967 1161 2001
rect 1161 1967 1195 2001
rect 1017 1929 1195 1967
rect 1017 1895 1051 1929
rect 1051 1895 1089 1929
rect 1089 1895 1123 1929
rect 1123 1895 1161 1929
rect 1161 1895 1195 1929
rect 1017 1857 1195 1895
rect 1017 1823 1051 1857
rect 1051 1823 1089 1857
rect 1089 1823 1123 1857
rect 1123 1823 1161 1857
rect 1161 1823 1195 1857
rect 1017 1785 1195 1823
rect 1017 1751 1051 1785
rect 1051 1751 1089 1785
rect 1089 1751 1123 1785
rect 1123 1751 1161 1785
rect 1161 1751 1195 1785
rect 1017 1713 1195 1751
rect 1017 1679 1051 1713
rect 1051 1679 1089 1713
rect 1089 1679 1123 1713
rect 1123 1679 1161 1713
rect 1161 1679 1195 1713
rect 1017 1641 1195 1679
rect 1017 1607 1051 1641
rect 1051 1607 1089 1641
rect 1089 1607 1123 1641
rect 1123 1607 1161 1641
rect 1161 1607 1195 1641
rect 1017 1569 1195 1607
rect 1017 1535 1051 1569
rect 1051 1535 1089 1569
rect 1089 1535 1123 1569
rect 1123 1535 1161 1569
rect 1161 1535 1195 1569
rect 1017 1497 1195 1535
rect 1017 1463 1051 1497
rect 1051 1463 1089 1497
rect 1089 1463 1123 1497
rect 1123 1463 1161 1497
rect 1161 1463 1195 1497
rect 1017 1425 1195 1463
rect 1017 1391 1051 1425
rect 1051 1391 1089 1425
rect 1089 1391 1123 1425
rect 1123 1391 1161 1425
rect 1161 1391 1195 1425
rect 1017 1353 1195 1391
rect 1017 1319 1051 1353
rect 1051 1319 1089 1353
rect 1089 1319 1123 1353
rect 1123 1319 1161 1353
rect 1161 1319 1195 1353
rect 1017 1281 1195 1319
rect 1017 1247 1051 1281
rect 1051 1247 1089 1281
rect 1089 1247 1123 1281
rect 1123 1247 1161 1281
rect 1161 1247 1195 1281
rect 1017 1209 1195 1247
rect 1017 1175 1051 1209
rect 1051 1175 1089 1209
rect 1089 1175 1123 1209
rect 1123 1175 1161 1209
rect 1161 1175 1195 1209
rect 1017 1137 1195 1175
rect 1017 1103 1051 1137
rect 1051 1103 1089 1137
rect 1089 1103 1123 1137
rect 1123 1103 1161 1137
rect 1161 1103 1195 1137
rect 1017 1065 1195 1103
rect 1017 1031 1051 1065
rect 1051 1031 1089 1065
rect 1089 1031 1123 1065
rect 1123 1031 1161 1065
rect 1161 1031 1195 1065
rect 1017 993 1195 1031
rect 1017 959 1051 993
rect 1051 959 1089 993
rect 1089 959 1123 993
rect 1123 959 1161 993
rect 1161 959 1195 993
rect 1017 921 1195 959
rect 1017 887 1051 921
rect 1051 887 1089 921
rect 1089 887 1123 921
rect 1123 887 1161 921
rect 1161 887 1195 921
rect 1017 849 1195 887
rect 1017 815 1051 849
rect 1051 815 1089 849
rect 1089 815 1123 849
rect 1123 815 1161 849
rect 1161 815 1195 849
rect 1017 777 1195 815
rect 1017 743 1051 777
rect 1051 743 1089 777
rect 1089 743 1123 777
rect 1123 743 1161 777
rect 1161 743 1195 777
rect 1017 705 1195 743
rect 1017 671 1051 705
rect 1051 671 1089 705
rect 1089 671 1123 705
rect 1123 671 1161 705
rect 1161 671 1195 705
rect 1017 633 1195 671
rect 1017 599 1051 633
rect 1051 599 1089 633
rect 1089 599 1123 633
rect 1123 599 1161 633
rect 1161 599 1195 633
rect 1017 561 1195 599
rect 1017 527 1051 561
rect 1051 527 1089 561
rect 1089 527 1123 561
rect 1123 527 1161 561
rect 1161 527 1195 561
rect 1017 489 1195 527
rect 1017 455 1051 489
rect 1051 455 1089 489
rect 1089 455 1123 489
rect 1123 455 1161 489
rect 1161 455 1195 489
rect 1017 417 1195 455
rect 1017 383 1051 417
rect 1051 383 1089 417
rect 1089 383 1123 417
rect 1123 383 1161 417
rect 1161 383 1195 417
rect 1017 345 1195 383
rect 1017 311 1051 345
rect 1051 311 1089 345
rect 1089 311 1123 345
rect 1123 311 1161 345
rect 1161 311 1195 345
rect 1017 273 1195 311
rect 1017 239 1051 273
rect 1051 239 1089 273
rect 1089 239 1123 273
rect 1123 239 1161 273
rect 1161 239 1195 273
rect 1017 201 1195 239
rect 1017 167 1051 201
rect 1051 167 1089 201
rect 1089 167 1123 201
rect 1123 167 1161 201
rect 1161 167 1195 201
rect 1017 129 1195 167
rect 1017 95 1051 129
rect 1051 95 1089 129
rect 1089 95 1123 129
rect 1123 95 1161 129
rect 1161 95 1195 129
rect 1017 57 1195 95
rect 1017 23 1051 57
rect 1051 23 1089 57
rect 1089 23 1123 57
rect 1123 23 1161 57
rect 1161 23 1195 57
<< metal1 >>
rect 215 8090 993 8096
rect 215 8056 227 8090
rect 261 8056 299 8090
rect 333 8056 371 8090
rect 405 8056 443 8090
rect 477 8056 515 8090
rect 549 8056 587 8090
rect 621 8056 659 8090
rect 693 8056 731 8090
rect 765 8056 803 8090
rect 837 8056 875 8090
rect 909 8056 947 8090
rect 981 8056 993 8090
rect 215 8050 993 8056
rect 7 7977 197 7989
rect 7 23 13 7977
rect 191 23 197 7977
rect 7 11 197 23
rect 1011 7977 1201 7989
rect 1011 23 1017 7977
rect 1195 23 1201 7977
rect 1011 11 1201 23
<< end >>
