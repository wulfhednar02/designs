magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< error_s >>
rect 1108 4544 1178 4572
rect 1362 4047 1432 4075
rect 1108 3550 1178 3578
rect 1362 3053 1432 3081
rect 1108 2556 1178 2584
rect 1362 2059 1432 2087
rect 1108 1562 1178 1590
rect 1362 1065 1432 1093
<< metal1 >>
rect 864 4603 914 5024
rect 1111 4970 1175 4976
rect 1111 4918 1117 4970
rect 1169 4918 1175 4970
rect 1111 4898 1175 4918
rect 1111 4846 1117 4898
rect 1169 4846 1175 4898
rect 1111 4826 1175 4846
rect 1111 4774 1117 4826
rect 1169 4774 1175 4826
rect 1111 4754 1175 4774
rect 1111 4702 1117 4754
rect 1169 4702 1175 4754
rect 1111 4682 1175 4702
rect 1111 4630 1117 4682
rect 1169 4630 1175 4682
rect 1111 4610 1175 4630
rect 1111 4558 1117 4610
rect 1169 4558 1175 4610
rect 1111 4552 1175 4558
rect 610 4106 660 4527
rect 864 4056 1422 4493
rect 356 3609 406 4030
rect 610 3559 1422 3996
rect 102 3112 152 3533
rect 356 3062 1422 3499
rect 102 2565 1422 3002
rect 102 2068 1422 2505
rect 102 1537 152 1958
rect 356 1571 1422 2008
rect 356 1040 406 1461
rect 610 1074 1422 1511
rect 610 543 660 964
rect 864 577 1422 1014
rect 864 46 914 467
rect 1111 463 1175 469
rect 1111 411 1117 463
rect 1169 411 1175 463
rect 1111 391 1175 411
rect 1111 339 1117 391
rect 1169 339 1175 391
rect 1111 319 1175 339
rect 1111 267 1117 319
rect 1169 267 1175 319
rect 1111 247 1175 267
rect 1111 195 1117 247
rect 1169 195 1175 247
rect 1111 175 1175 195
rect 1111 123 1117 175
rect 1169 123 1175 175
rect 1111 103 1175 123
rect 1111 51 1117 103
rect 1169 51 1175 103
rect 1111 45 1175 51
<< via1 >>
rect 1117 4918 1169 4970
rect 1117 4846 1169 4898
rect 1117 4774 1169 4826
rect 1117 4702 1169 4754
rect 1117 4630 1169 4682
rect 1117 4558 1169 4610
rect 1117 411 1169 463
rect 1117 339 1169 391
rect 1117 267 1169 319
rect 1117 195 1169 247
rect 1117 123 1169 175
rect 1117 51 1169 103
<< metal2 >>
rect 1111 4970 1175 4976
rect 1111 4918 1117 4970
rect 1169 4918 1175 4970
rect 1111 4898 1175 4918
rect 1111 4846 1117 4898
rect 1169 4846 1175 4898
rect 1111 4826 1175 4846
rect 1111 4774 1117 4826
rect 1169 4774 1175 4826
rect 1111 4754 1175 4774
rect 1111 4702 1117 4754
rect 1169 4702 1175 4754
rect 1111 4682 1175 4702
rect 1111 4630 1117 4682
rect 1169 4630 1175 4682
rect 1111 4610 1175 4630
rect 1111 4558 1117 4610
rect 1169 4558 1175 4610
rect 1111 4552 1175 4558
rect 1111 463 1175 469
rect 1111 411 1117 463
rect 1169 411 1175 463
rect 1111 391 1175 411
rect 1111 339 1117 391
rect 1169 339 1175 391
rect 1111 319 1175 339
rect 1111 267 1117 319
rect 1169 267 1175 319
rect 1111 247 1175 267
rect 1111 195 1117 247
rect 1169 195 1175 247
rect 1111 175 1175 195
rect 1111 123 1117 175
rect 1169 123 1175 175
rect 1111 103 1175 123
rect 1111 51 1117 103
rect 1169 51 1175 103
rect 1111 45 1175 51
use res_poly$5  res_poly$5_0
timestamp 1698982078
transform 1 0 508 0 1 497
box 92 40 162 1004
use res_poly$5  res_poly$5_1
timestamp 1698982078
transform 1 0 762 0 1 0
box 92 40 162 1004
use res_poly$5  res_poly$5_2
timestamp 1698982078
transform 1 0 508 0 1 3529
box 92 40 162 1004
use res_poly$5  res_poly$5_3
timestamp 1698982078
transform 1 0 762 0 1 4026
box 92 40 162 1004
use res_poly$5  res_poly$5_4
timestamp 1698982078
transform 1 0 1016 0 1 0
box 92 40 162 1004
use res_poly$5  res_poly$5_5
timestamp 1698982078
transform 1 0 0 0 1 1491
box 92 40 162 1004
use res_poly$5  res_poly$5_6
timestamp 1698982078
transform 1 0 254 0 1 3032
box 92 40 162 1004
use res_poly$5  res_poly$5_7
timestamp 1698982078
transform 1 0 254 0 1 994
box 92 40 162 1004
use res_poly$5  res_poly$5_8
timestamp 1698982078
transform 1 0 0 0 1 2535
box 92 40 162 1004
use res_poly  res_poly_0
timestamp 1698982078
transform 1 0 1270 0 1 1541
box 92 40 162 954
use res_poly  res_poly_1
timestamp 1698982078
transform 1 0 1016 0 1 4026
box 92 40 162 954
use res_poly  res_poly_2
timestamp 1698982078
transform 1 0 1016 0 1 3032
box 92 40 162 954
use res_poly  res_poly_3
timestamp 1698982078
transform 1 0 1270 0 1 3529
box 92 40 162 954
use res_poly  res_poly_4
timestamp 1698982078
transform 1 0 1270 0 1 2535
box 92 40 162 954
use res_poly  res_poly_5
timestamp 1698982078
transform 1 0 1270 0 1 547
box 92 40 162 954
use res_poly  res_poly_6
timestamp 1698982078
transform 1 0 1016 0 1 1044
box 92 40 162 954
use res_poly  res_poly_7
timestamp 1698982078
transform 1 0 1016 0 1 2038
box 92 40 162 954
<< labels >>
flabel metal1 s 864 4056 1422 4492 0 FreeSans 44 0 0 0 OUT
port 2 nsew
flabel metal1 s 1007 4278 1007 4278 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 993 4467 993 4467 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 356 3609 406 4030 0 FreeSans 44 0 0 0 DAC5
port 3 nsew
flabel metal1 s 381 3822 381 3822 0 FreeSans 44 0 0 0 DAC5
flabel metal1 s 378 4002 378 4002 0 FreeSans 44 0 0 0 DAC5
flabel metal1 s 610 4106 660 4527 0 FreeSans 44 0 0 0 DAC6
port 4 nsew
flabel metal1 s 864 4603 914 5024 0 FreeSans 44 0 0 0 DAC7
port 5 nsew
flabel metal1 s 633 4499 633 4499 0 FreeSans 44 0 0 0 DAC6
flabel metal1 s 635 4314 635 4314 0 FreeSans 44 0 0 0 DAC6
flabel metal1 s 887 4633 887 4633 0 FreeSans 44 0 0 0 DAC7
flabel metal1 s 887 4814 887 4814 0 FreeSans 44 0 0 0 DAC7
flabel metal1 s 1266 4456 1266 4456 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 1265 4291 1265 4291 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 1266 4098 1266 4098 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 102 3112 152 3533 0 FreeSans 44 0 0 0 DAC4
port 6 nsew
flabel metal1 s 125 3322 125 3322 0 FreeSans 44 0 0 0 DAC4
flabel metal1 s 125 3142 125 3142 0 FreeSans 44 0 0 0 DAC4
flabel metal1 s 102 1537 152 1957 0 FreeSans 44 0 0 0 DAC3
port 7 nsew
flabel metal1 s 128 1753 128 1753 0 FreeSans 44 0 0 0 DAC3
flabel metal1 s 126 1568 126 1568 0 FreeSans 44 0 0 0 DAC3
flabel metal1 s 356 1040 406 1460 0 FreeSans 44 0 0 0 DAC2
port 8 nsew
flabel metal1 s 379 1429 379 1429 0 FreeSans 44 0 0 0 DAC2
flabel metal1 s 382 1072 382 1072 0 FreeSans 44 0 0 0 DAC2
flabel metal1 s 610 543 660 963 0 FreeSans 44 0 0 0 DAC1
port 9 nsew
flabel metal1 s 638 937 638 937 0 FreeSans 44 0 0 0 DAC1
flabel metal1 s 636 574 636 574 0 FreeSans 44 0 0 0 DAC1
flabel metal1 s 864 46 914 466 0 FreeSans 44 0 0 0 DAC0
port 10 nsew
flabel metal1 s 888 437 888 437 0 FreeSans 44 0 0 0 DAC0
flabel metal1 s 888 77 888 77 0 FreeSans 44 0 0 0 DAC0
flabel metal2 s 1111 4552 1175 4976 0 FreeSans 44 0 0 0 VDD
port 12 nsew
flabel metal2 s 1142 4767 1142 4767 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 1142 4583 1142 4583 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 1111 45 1175 469 0 FreeSans 44 0 0 0 VSS
port 13 nsew
flabel metal2 s 1140 75 1140 75 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 1141 436 1141 436 0 FreeSans 44 0 0 0 VSS
<< end >>
