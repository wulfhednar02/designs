magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< nwell >>
rect 0 309 2100 630
<< pwell >>
rect 39 69 1989 251
rect 68 31 102 69
<< scnmos >>
rect 117 95 147 225
rect 201 95 231 225
rect 285 95 315 225
rect 369 95 399 225
rect 453 95 483 225
rect 537 95 567 225
rect 621 95 651 225
rect 705 95 735 225
rect 789 95 819 225
rect 873 95 903 225
rect 957 95 987 225
rect 1041 95 1071 225
rect 1125 95 1155 225
rect 1209 95 1239 225
rect 1293 95 1323 225
rect 1377 95 1407 225
rect 1461 95 1491 225
rect 1545 95 1575 225
rect 1629 95 1659 225
rect 1713 95 1743 225
rect 1797 95 1827 225
rect 1881 95 1911 225
<< scpmoshvt >>
rect 117 345 147 545
rect 201 345 231 545
rect 285 345 315 545
rect 369 345 399 545
rect 453 345 483 545
rect 537 345 567 545
rect 621 345 651 545
rect 705 345 735 545
rect 789 345 819 545
rect 873 345 903 545
rect 957 345 987 545
rect 1041 345 1071 545
rect 1125 345 1155 545
rect 1209 345 1239 545
rect 1293 345 1323 545
rect 1377 345 1407 545
rect 1461 345 1491 545
rect 1545 345 1575 545
rect 1629 345 1659 545
rect 1713 345 1743 545
rect 1797 345 1827 545
rect 1881 345 1911 545
<< ndiff >>
rect 65 213 117 225
rect 65 179 73 213
rect 107 179 117 213
rect 65 145 117 179
rect 65 111 73 145
rect 107 111 117 145
rect 65 95 117 111
rect 147 213 201 225
rect 147 179 157 213
rect 191 179 201 213
rect 147 145 201 179
rect 147 111 157 145
rect 191 111 201 145
rect 147 95 201 111
rect 231 145 285 225
rect 231 111 241 145
rect 275 111 285 145
rect 231 95 285 111
rect 315 213 369 225
rect 315 179 325 213
rect 359 179 369 213
rect 315 145 369 179
rect 315 111 325 145
rect 359 111 369 145
rect 315 95 369 111
rect 399 145 453 225
rect 399 111 409 145
rect 443 111 453 145
rect 399 95 453 111
rect 483 213 537 225
rect 483 179 493 213
rect 527 179 537 213
rect 483 145 537 179
rect 483 111 493 145
rect 527 111 537 145
rect 483 95 537 111
rect 567 145 621 225
rect 567 111 577 145
rect 611 111 621 145
rect 567 95 621 111
rect 651 213 705 225
rect 651 179 661 213
rect 695 179 705 213
rect 651 145 705 179
rect 651 111 661 145
rect 695 111 705 145
rect 651 95 705 111
rect 735 145 789 225
rect 735 111 745 145
rect 779 111 789 145
rect 735 95 789 111
rect 819 213 873 225
rect 819 179 829 213
rect 863 179 873 213
rect 819 145 873 179
rect 819 111 829 145
rect 863 111 873 145
rect 819 95 873 111
rect 903 145 957 225
rect 903 111 913 145
rect 947 111 957 145
rect 903 95 957 111
rect 987 213 1041 225
rect 987 179 997 213
rect 1031 179 1041 213
rect 987 145 1041 179
rect 987 111 997 145
rect 1031 111 1041 145
rect 987 95 1041 111
rect 1071 145 1125 225
rect 1071 111 1081 145
rect 1115 111 1125 145
rect 1071 95 1125 111
rect 1155 213 1209 225
rect 1155 179 1165 213
rect 1199 179 1209 213
rect 1155 145 1209 179
rect 1155 111 1165 145
rect 1199 111 1209 145
rect 1155 95 1209 111
rect 1239 145 1293 225
rect 1239 111 1249 145
rect 1283 111 1293 145
rect 1239 95 1293 111
rect 1323 213 1377 225
rect 1323 179 1333 213
rect 1367 179 1377 213
rect 1323 145 1377 179
rect 1323 111 1333 145
rect 1367 111 1377 145
rect 1323 95 1377 111
rect 1407 145 1461 225
rect 1407 111 1417 145
rect 1451 111 1461 145
rect 1407 95 1461 111
rect 1491 213 1545 225
rect 1491 179 1501 213
rect 1535 179 1545 213
rect 1491 145 1545 179
rect 1491 111 1501 145
rect 1535 111 1545 145
rect 1491 95 1545 111
rect 1575 145 1629 225
rect 1575 111 1585 145
rect 1619 111 1629 145
rect 1575 95 1629 111
rect 1659 213 1713 225
rect 1659 179 1669 213
rect 1703 179 1713 213
rect 1659 145 1713 179
rect 1659 111 1669 145
rect 1703 111 1713 145
rect 1659 95 1713 111
rect 1743 145 1797 225
rect 1743 111 1753 145
rect 1787 111 1797 145
rect 1743 95 1797 111
rect 1827 213 1881 225
rect 1827 179 1837 213
rect 1871 179 1881 213
rect 1827 145 1881 179
rect 1827 111 1837 145
rect 1871 111 1881 145
rect 1827 95 1881 111
rect 1911 145 1963 225
rect 1911 111 1921 145
rect 1955 111 1963 145
rect 1911 95 1963 111
<< pdiff >>
rect 65 533 117 545
rect 65 499 73 533
rect 107 499 117 533
rect 65 465 117 499
rect 65 431 73 465
rect 107 431 117 465
rect 65 397 117 431
rect 65 363 73 397
rect 107 363 117 397
rect 65 345 117 363
rect 147 527 201 545
rect 147 493 157 527
rect 191 493 201 527
rect 147 459 201 493
rect 147 425 157 459
rect 191 425 201 459
rect 147 391 201 425
rect 147 357 157 391
rect 191 357 201 391
rect 147 345 201 357
rect 231 533 285 545
rect 231 499 241 533
rect 275 499 285 533
rect 231 465 285 499
rect 231 431 241 465
rect 275 431 285 465
rect 231 345 285 431
rect 315 527 369 545
rect 315 493 325 527
rect 359 493 369 527
rect 315 459 369 493
rect 315 425 325 459
rect 359 425 369 459
rect 315 391 369 425
rect 315 357 325 391
rect 359 357 369 391
rect 315 345 369 357
rect 399 533 453 545
rect 399 499 409 533
rect 443 499 453 533
rect 399 465 453 499
rect 399 431 409 465
rect 443 431 453 465
rect 399 345 453 431
rect 483 527 537 545
rect 483 493 493 527
rect 527 493 537 527
rect 483 459 537 493
rect 483 425 493 459
rect 527 425 537 459
rect 483 391 537 425
rect 483 357 493 391
rect 527 357 537 391
rect 483 345 537 357
rect 567 533 621 545
rect 567 499 577 533
rect 611 499 621 533
rect 567 465 621 499
rect 567 431 577 465
rect 611 431 621 465
rect 567 345 621 431
rect 651 527 705 545
rect 651 493 661 527
rect 695 493 705 527
rect 651 459 705 493
rect 651 425 661 459
rect 695 425 705 459
rect 651 391 705 425
rect 651 357 661 391
rect 695 357 705 391
rect 651 345 705 357
rect 735 533 789 545
rect 735 499 745 533
rect 779 499 789 533
rect 735 465 789 499
rect 735 431 745 465
rect 779 431 789 465
rect 735 345 789 431
rect 819 527 873 545
rect 819 493 829 527
rect 863 493 873 527
rect 819 459 873 493
rect 819 425 829 459
rect 863 425 873 459
rect 819 391 873 425
rect 819 357 829 391
rect 863 357 873 391
rect 819 345 873 357
rect 903 533 957 545
rect 903 499 913 533
rect 947 499 957 533
rect 903 465 957 499
rect 903 431 913 465
rect 947 431 957 465
rect 903 345 957 431
rect 987 527 1041 545
rect 987 493 997 527
rect 1031 493 1041 527
rect 987 459 1041 493
rect 987 425 997 459
rect 1031 425 1041 459
rect 987 391 1041 425
rect 987 357 997 391
rect 1031 357 1041 391
rect 987 345 1041 357
rect 1071 533 1125 545
rect 1071 499 1081 533
rect 1115 499 1125 533
rect 1071 465 1125 499
rect 1071 431 1081 465
rect 1115 431 1125 465
rect 1071 345 1125 431
rect 1155 527 1209 545
rect 1155 493 1165 527
rect 1199 493 1209 527
rect 1155 459 1209 493
rect 1155 425 1165 459
rect 1199 425 1209 459
rect 1155 391 1209 425
rect 1155 357 1165 391
rect 1199 357 1209 391
rect 1155 345 1209 357
rect 1239 533 1293 545
rect 1239 499 1249 533
rect 1283 499 1293 533
rect 1239 465 1293 499
rect 1239 431 1249 465
rect 1283 431 1293 465
rect 1239 345 1293 431
rect 1323 527 1377 545
rect 1323 493 1333 527
rect 1367 493 1377 527
rect 1323 459 1377 493
rect 1323 425 1333 459
rect 1367 425 1377 459
rect 1323 391 1377 425
rect 1323 357 1333 391
rect 1367 357 1377 391
rect 1323 345 1377 357
rect 1407 533 1461 545
rect 1407 499 1417 533
rect 1451 499 1461 533
rect 1407 465 1461 499
rect 1407 431 1417 465
rect 1451 431 1461 465
rect 1407 345 1461 431
rect 1491 527 1545 545
rect 1491 493 1501 527
rect 1535 493 1545 527
rect 1491 459 1545 493
rect 1491 425 1501 459
rect 1535 425 1545 459
rect 1491 391 1545 425
rect 1491 357 1501 391
rect 1535 357 1545 391
rect 1491 345 1545 357
rect 1575 533 1629 545
rect 1575 499 1585 533
rect 1619 499 1629 533
rect 1575 465 1629 499
rect 1575 431 1585 465
rect 1619 431 1629 465
rect 1575 345 1629 431
rect 1659 527 1713 545
rect 1659 493 1669 527
rect 1703 493 1713 527
rect 1659 459 1713 493
rect 1659 425 1669 459
rect 1703 425 1713 459
rect 1659 391 1713 425
rect 1659 357 1669 391
rect 1703 357 1713 391
rect 1659 345 1713 357
rect 1743 533 1797 545
rect 1743 499 1753 533
rect 1787 499 1797 533
rect 1743 465 1797 499
rect 1743 431 1753 465
rect 1787 431 1797 465
rect 1743 345 1797 431
rect 1827 527 1881 545
rect 1827 493 1837 527
rect 1871 493 1881 527
rect 1827 459 1881 493
rect 1827 425 1837 459
rect 1871 425 1881 459
rect 1827 391 1881 425
rect 1827 357 1837 391
rect 1871 357 1881 391
rect 1827 345 1881 357
rect 1911 533 1963 545
rect 1911 499 1921 533
rect 1955 499 1963 533
rect 1911 465 1963 499
rect 1911 431 1921 465
rect 1955 431 1963 465
rect 1911 345 1963 431
<< ndiffc >>
rect 73 179 107 213
rect 73 111 107 145
rect 157 179 191 213
rect 157 111 191 145
rect 241 111 275 145
rect 325 179 359 213
rect 325 111 359 145
rect 409 111 443 145
rect 493 179 527 213
rect 493 111 527 145
rect 577 111 611 145
rect 661 179 695 213
rect 661 111 695 145
rect 745 111 779 145
rect 829 179 863 213
rect 829 111 863 145
rect 913 111 947 145
rect 997 179 1031 213
rect 997 111 1031 145
rect 1081 111 1115 145
rect 1165 179 1199 213
rect 1165 111 1199 145
rect 1249 111 1283 145
rect 1333 179 1367 213
rect 1333 111 1367 145
rect 1417 111 1451 145
rect 1501 179 1535 213
rect 1501 111 1535 145
rect 1585 111 1619 145
rect 1669 179 1703 213
rect 1669 111 1703 145
rect 1753 111 1787 145
rect 1837 179 1871 213
rect 1837 111 1871 145
rect 1921 111 1955 145
<< pdiffc >>
rect 73 499 107 533
rect 73 431 107 465
rect 73 363 107 397
rect 157 493 191 527
rect 157 425 191 459
rect 157 357 191 391
rect 241 499 275 533
rect 241 431 275 465
rect 325 493 359 527
rect 325 425 359 459
rect 325 357 359 391
rect 409 499 443 533
rect 409 431 443 465
rect 493 493 527 527
rect 493 425 527 459
rect 493 357 527 391
rect 577 499 611 533
rect 577 431 611 465
rect 661 493 695 527
rect 661 425 695 459
rect 661 357 695 391
rect 745 499 779 533
rect 745 431 779 465
rect 829 493 863 527
rect 829 425 863 459
rect 829 357 863 391
rect 913 499 947 533
rect 913 431 947 465
rect 997 493 1031 527
rect 997 425 1031 459
rect 997 357 1031 391
rect 1081 499 1115 533
rect 1081 431 1115 465
rect 1165 493 1199 527
rect 1165 425 1199 459
rect 1165 357 1199 391
rect 1249 499 1283 533
rect 1249 431 1283 465
rect 1333 493 1367 527
rect 1333 425 1367 459
rect 1333 357 1367 391
rect 1417 499 1451 533
rect 1417 431 1451 465
rect 1501 493 1535 527
rect 1501 425 1535 459
rect 1501 357 1535 391
rect 1585 499 1619 533
rect 1585 431 1619 465
rect 1669 493 1703 527
rect 1669 425 1703 459
rect 1669 357 1703 391
rect 1753 499 1787 533
rect 1753 431 1787 465
rect 1837 493 1871 527
rect 1837 425 1871 459
rect 1837 357 1871 391
rect 1921 499 1955 533
rect 1921 431 1955 465
<< poly >>
rect 117 545 147 571
rect 201 545 231 571
rect 285 545 315 571
rect 369 545 399 571
rect 453 545 483 571
rect 537 545 567 571
rect 621 545 651 571
rect 705 545 735 571
rect 789 545 819 571
rect 873 545 903 571
rect 957 545 987 571
rect 1041 545 1071 571
rect 1125 545 1155 571
rect 1209 545 1239 571
rect 1293 545 1323 571
rect 1377 545 1407 571
rect 1461 545 1491 571
rect 1545 545 1575 571
rect 1629 545 1659 571
rect 1713 545 1743 571
rect 1797 545 1827 571
rect 1881 545 1911 571
rect 117 307 147 345
rect 201 307 231 345
rect 285 307 315 345
rect 369 307 399 345
rect 453 307 483 345
rect 537 307 567 345
rect 117 297 567 307
rect 117 263 141 297
rect 175 263 209 297
rect 243 263 277 297
rect 311 263 345 297
rect 379 263 413 297
rect 447 263 481 297
rect 515 263 567 297
rect 117 253 567 263
rect 117 225 147 253
rect 201 225 231 253
rect 285 225 315 253
rect 369 225 399 253
rect 453 225 483 253
rect 537 225 567 253
rect 621 307 651 345
rect 705 307 735 345
rect 789 307 819 345
rect 873 307 903 345
rect 957 307 987 345
rect 1041 307 1071 345
rect 1125 307 1155 345
rect 1209 307 1239 345
rect 1293 307 1323 345
rect 1377 307 1407 345
rect 1461 307 1491 345
rect 1545 307 1575 345
rect 1629 307 1659 345
rect 1713 307 1743 345
rect 1797 307 1827 345
rect 1881 307 1911 345
rect 621 297 1915 307
rect 621 263 641 297
rect 675 263 709 297
rect 743 263 777 297
rect 811 263 845 297
rect 879 263 913 297
rect 947 263 981 297
rect 1015 263 1049 297
rect 1083 263 1117 297
rect 1151 263 1185 297
rect 1219 263 1253 297
rect 1287 263 1321 297
rect 1355 263 1389 297
rect 1423 263 1457 297
rect 1491 263 1525 297
rect 1559 263 1593 297
rect 1627 263 1661 297
rect 1695 263 1729 297
rect 1763 263 1797 297
rect 1831 263 1865 297
rect 1899 263 1915 297
rect 621 253 1915 263
rect 621 225 651 253
rect 705 225 735 253
rect 789 225 819 253
rect 873 225 903 253
rect 957 225 987 253
rect 1041 225 1071 253
rect 1125 225 1155 253
rect 1209 225 1239 253
rect 1293 225 1323 253
rect 1377 225 1407 253
rect 1461 225 1491 253
rect 1545 225 1575 253
rect 1629 225 1659 253
rect 1713 225 1743 253
rect 1797 225 1827 253
rect 1881 225 1911 253
rect 117 69 147 95
rect 201 69 231 95
rect 285 69 315 95
rect 369 69 399 95
rect 453 69 483 95
rect 537 69 567 95
rect 621 69 651 95
rect 705 69 735 95
rect 789 69 819 95
rect 873 69 903 95
rect 957 69 987 95
rect 1041 69 1071 95
rect 1125 69 1155 95
rect 1209 69 1239 95
rect 1293 69 1323 95
rect 1377 69 1407 95
rect 1461 69 1491 95
rect 1545 69 1575 95
rect 1629 69 1659 95
rect 1713 69 1743 95
rect 1797 69 1827 95
rect 1881 69 1911 95
<< polycont >>
rect 141 263 175 297
rect 209 263 243 297
rect 277 263 311 297
rect 345 263 379 297
rect 413 263 447 297
rect 481 263 515 297
rect 641 263 675 297
rect 709 263 743 297
rect 777 263 811 297
rect 845 263 879 297
rect 913 263 947 297
rect 981 263 1015 297
rect 1049 263 1083 297
rect 1117 263 1151 297
rect 1185 263 1219 297
rect 1253 263 1287 297
rect 1321 263 1355 297
rect 1389 263 1423 297
rect 1457 263 1491 297
rect 1525 263 1559 297
rect 1593 263 1627 297
rect 1661 263 1695 297
rect 1729 263 1763 297
rect 1797 263 1831 297
rect 1865 263 1899 297
<< locali >>
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 343 609
rect 377 575 435 609
rect 469 575 527 609
rect 561 575 619 609
rect 653 575 711 609
rect 745 575 803 609
rect 837 575 895 609
rect 929 575 987 609
rect 1021 575 1079 609
rect 1113 575 1171 609
rect 1205 575 1263 609
rect 1297 575 1355 609
rect 1389 575 1447 609
rect 1481 575 1539 609
rect 1573 575 1631 609
rect 1665 575 1723 609
rect 1757 575 1815 609
rect 1849 575 1907 609
rect 1941 575 1999 609
rect 2033 575 2062 609
rect 73 533 107 575
rect 73 465 107 499
rect 73 397 107 431
rect 73 337 107 363
rect 141 527 207 541
rect 141 493 157 527
rect 191 493 207 527
rect 141 459 207 493
rect 141 425 157 459
rect 191 425 207 459
rect 141 391 207 425
rect 241 533 275 575
rect 241 465 275 499
rect 241 415 275 431
rect 309 527 375 541
rect 309 493 325 527
rect 359 493 375 527
rect 309 459 375 493
rect 309 425 325 459
rect 359 425 375 459
rect 141 357 157 391
rect 191 371 207 391
rect 309 391 375 425
rect 409 533 443 575
rect 409 465 443 499
rect 409 415 443 431
rect 477 527 543 541
rect 477 493 493 527
rect 527 493 543 527
rect 477 459 543 493
rect 477 425 493 459
rect 527 425 543 459
rect 309 371 325 391
rect 191 357 325 371
rect 359 371 375 391
rect 477 391 543 425
rect 577 533 611 575
rect 577 465 611 499
rect 577 415 611 431
rect 645 527 711 541
rect 645 493 661 527
rect 695 493 711 527
rect 645 459 711 493
rect 645 425 661 459
rect 695 425 711 459
rect 477 371 493 391
rect 359 357 493 371
rect 527 371 543 391
rect 645 391 711 425
rect 745 533 779 575
rect 745 465 779 499
rect 745 415 779 431
rect 813 527 879 541
rect 813 493 829 527
rect 863 493 879 527
rect 813 459 879 493
rect 813 425 829 459
rect 863 425 879 459
rect 527 357 611 371
rect 141 337 611 357
rect 645 357 661 391
rect 695 371 711 391
rect 813 391 879 425
rect 913 533 947 575
rect 913 465 947 499
rect 913 415 947 431
rect 981 527 1047 541
rect 981 493 997 527
rect 1031 493 1047 527
rect 981 459 1047 493
rect 981 425 997 459
rect 1031 425 1047 459
rect 813 371 829 391
rect 695 357 829 371
rect 863 371 879 391
rect 981 391 1047 425
rect 1081 533 1115 575
rect 1081 465 1115 499
rect 1081 415 1115 431
rect 1149 527 1215 541
rect 1149 493 1165 527
rect 1199 493 1215 527
rect 1149 459 1215 493
rect 1149 425 1165 459
rect 1199 425 1215 459
rect 981 371 997 391
rect 863 357 997 371
rect 1031 371 1047 391
rect 1149 391 1215 425
rect 1249 533 1283 575
rect 1249 465 1283 499
rect 1249 415 1283 431
rect 1317 527 1383 541
rect 1317 493 1333 527
rect 1367 493 1383 527
rect 1317 459 1383 493
rect 1317 425 1333 459
rect 1367 425 1383 459
rect 1149 371 1165 391
rect 1031 357 1165 371
rect 1199 371 1215 391
rect 1317 391 1383 425
rect 1417 533 1451 575
rect 1417 465 1451 499
rect 1417 415 1451 431
rect 1485 527 1551 541
rect 1485 493 1501 527
rect 1535 493 1551 527
rect 1485 459 1551 493
rect 1485 425 1501 459
rect 1535 425 1551 459
rect 1317 371 1333 391
rect 1199 357 1333 371
rect 1367 371 1383 391
rect 1485 391 1551 425
rect 1585 533 1619 575
rect 1585 465 1619 499
rect 1585 415 1619 431
rect 1653 527 1719 541
rect 1653 493 1669 527
rect 1703 493 1719 527
rect 1653 459 1719 493
rect 1653 425 1669 459
rect 1703 425 1719 459
rect 1485 371 1501 391
rect 1367 357 1501 371
rect 1535 371 1551 391
rect 1653 391 1719 425
rect 1753 533 1787 575
rect 1753 465 1787 499
rect 1753 415 1787 431
rect 1821 527 1887 541
rect 1821 493 1837 527
rect 1871 493 1887 527
rect 1821 459 1887 493
rect 1821 425 1837 459
rect 1871 425 1887 459
rect 1653 371 1669 391
rect 1535 357 1669 371
rect 1703 371 1719 391
rect 1821 391 1887 425
rect 1921 533 1955 575
rect 1921 465 1955 499
rect 1921 415 1955 431
rect 1821 371 1837 391
rect 1703 357 1837 371
rect 1871 371 1887 391
rect 1990 371 2045 520
rect 1871 357 2045 371
rect 645 337 2045 357
rect 576 303 611 337
rect 55 297 535 303
rect 55 263 141 297
rect 175 263 209 297
rect 243 263 277 297
rect 311 263 345 297
rect 379 263 413 297
rect 447 263 481 297
rect 515 263 535 297
rect 576 297 1920 303
rect 576 263 641 297
rect 675 263 709 297
rect 743 263 777 297
rect 811 263 845 297
rect 879 263 913 297
rect 947 263 981 297
rect 1015 263 1049 297
rect 1083 263 1117 297
rect 1151 263 1185 297
rect 1219 263 1253 297
rect 1287 263 1321 297
rect 1355 263 1389 297
rect 1423 263 1457 297
rect 1491 263 1525 297
rect 1559 263 1593 297
rect 1627 263 1661 297
rect 1695 263 1729 297
rect 1763 263 1797 297
rect 1831 263 1865 297
rect 1899 263 1920 297
rect 576 229 611 263
rect 1969 229 2045 337
rect 73 213 107 229
rect 73 145 107 179
rect 73 65 107 111
rect 141 213 611 229
rect 141 179 157 213
rect 191 195 325 213
rect 191 179 207 195
rect 141 145 207 179
rect 309 179 325 195
rect 359 195 493 213
rect 359 179 375 195
rect 141 111 157 145
rect 191 111 207 145
rect 141 100 207 111
rect 241 145 275 161
rect 241 65 275 111
rect 309 145 375 179
rect 477 179 493 195
rect 527 195 611 213
rect 645 213 2045 229
rect 527 179 543 195
rect 309 111 325 145
rect 359 111 375 145
rect 309 100 375 111
rect 409 145 443 161
rect 409 65 443 111
rect 477 145 543 179
rect 645 179 661 213
rect 695 195 829 213
rect 695 179 711 195
rect 477 111 493 145
rect 527 111 543 145
rect 477 100 543 111
rect 577 145 611 161
rect 577 65 611 111
rect 645 145 711 179
rect 813 179 829 195
rect 863 195 997 213
rect 863 179 879 195
rect 645 111 661 145
rect 695 111 711 145
rect 645 100 711 111
rect 745 145 779 161
rect 645 99 695 100
rect 745 65 779 111
rect 813 145 879 179
rect 981 179 997 195
rect 1031 195 1165 213
rect 1031 179 1047 195
rect 813 111 829 145
rect 863 111 879 145
rect 813 100 879 111
rect 913 145 947 161
rect 829 99 863 100
rect 913 65 947 111
rect 981 145 1047 179
rect 1149 179 1165 195
rect 1199 195 1333 213
rect 1199 179 1215 195
rect 981 111 997 145
rect 1031 111 1047 145
rect 981 100 1047 111
rect 1081 145 1115 161
rect 997 99 1031 100
rect 1081 65 1115 111
rect 1149 145 1215 179
rect 1317 179 1333 195
rect 1367 195 1501 213
rect 1367 179 1383 195
rect 1149 111 1165 145
rect 1199 111 1215 145
rect 1149 100 1215 111
rect 1249 145 1283 161
rect 1249 65 1283 111
rect 1317 145 1383 179
rect 1485 179 1501 195
rect 1535 195 1669 213
rect 1535 179 1551 195
rect 1317 111 1333 145
rect 1367 111 1383 145
rect 1317 100 1383 111
rect 1417 145 1451 161
rect 1417 65 1451 111
rect 1485 145 1551 179
rect 1653 179 1669 195
rect 1703 195 1837 213
rect 1703 179 1719 195
rect 1485 111 1501 145
rect 1535 111 1551 145
rect 1485 100 1551 111
rect 1585 145 1619 161
rect 1585 65 1619 111
rect 1653 145 1719 179
rect 1821 179 1837 195
rect 1871 195 2045 213
rect 1871 179 1887 195
rect 1653 111 1669 145
rect 1703 111 1719 145
rect 1653 100 1719 111
rect 1753 145 1787 161
rect 1753 65 1787 111
rect 1821 145 1887 179
rect 1821 111 1837 145
rect 1871 111 1887 145
rect 1821 100 1887 111
rect 1921 145 1955 161
rect 1990 121 2045 195
rect 1921 65 1955 111
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 343 65
rect 377 31 435 65
rect 469 31 527 65
rect 561 31 619 65
rect 653 31 711 65
rect 745 31 803 65
rect 837 31 895 65
rect 929 31 987 65
rect 1021 31 1079 65
rect 1113 31 1171 65
rect 1205 31 1263 65
rect 1297 31 1355 65
rect 1389 31 1447 65
rect 1481 31 1539 65
rect 1573 31 1631 65
rect 1665 31 1723 65
rect 1757 31 1815 65
rect 1849 31 1907 65
rect 1941 31 1999 65
rect 2033 31 2062 65
<< viali >>
rect 67 575 101 609
rect 159 575 193 609
rect 251 575 285 609
rect 343 575 377 609
rect 435 575 469 609
rect 527 575 561 609
rect 619 575 653 609
rect 711 575 745 609
rect 803 575 837 609
rect 895 575 929 609
rect 987 575 1021 609
rect 1079 575 1113 609
rect 1171 575 1205 609
rect 1263 575 1297 609
rect 1355 575 1389 609
rect 1447 575 1481 609
rect 1539 575 1573 609
rect 1631 575 1665 609
rect 1723 575 1757 609
rect 1815 575 1849 609
rect 1907 575 1941 609
rect 1999 575 2033 609
rect 67 31 101 65
rect 159 31 193 65
rect 251 31 285 65
rect 343 31 377 65
rect 435 31 469 65
rect 527 31 561 65
rect 619 31 653 65
rect 711 31 745 65
rect 803 31 837 65
rect 895 31 929 65
rect 987 31 1021 65
rect 1079 31 1113 65
rect 1171 31 1205 65
rect 1263 31 1297 65
rect 1355 31 1389 65
rect 1447 31 1481 65
rect 1539 31 1573 65
rect 1631 31 1665 65
rect 1723 31 1757 65
rect 1815 31 1849 65
rect 1907 31 1941 65
rect 1999 31 2033 65
<< metal1 >>
rect 38 609 2062 640
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 343 609
rect 377 575 435 609
rect 469 575 527 609
rect 561 575 619 609
rect 653 575 711 609
rect 745 575 803 609
rect 837 575 895 609
rect 929 575 987 609
rect 1021 575 1079 609
rect 1113 575 1171 609
rect 1205 575 1263 609
rect 1297 575 1355 609
rect 1389 575 1447 609
rect 1481 575 1539 609
rect 1573 575 1631 609
rect 1665 575 1723 609
rect 1757 575 1815 609
rect 1849 575 1907 609
rect 1941 575 1999 609
rect 2033 575 2062 609
rect 38 544 2062 575
rect 38 65 2062 96
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 343 65
rect 377 31 435 65
rect 469 31 527 65
rect 561 31 619 65
rect 653 31 711 65
rect 745 31 803 65
rect 837 31 895 65
rect 929 31 987 65
rect 1021 31 1079 65
rect 1113 31 1171 65
rect 1205 31 1263 65
rect 1297 31 1355 65
rect 1389 31 1447 65
rect 1481 31 1539 65
rect 1573 31 1631 65
rect 1665 31 1723 65
rect 1757 31 1815 65
rect 1849 31 1907 65
rect 1941 31 1999 65
rect 2033 31 2062 65
rect 38 0 2062 31
<< labels >>
flabel locali s 436 269 470 303 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel locali s 344 269 378 303 0 FreeSans 200 0 0 0 A
port 6 nsew
flabel locali s 1999 269 2033 303 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel locali s 1999 337 2033 371 0 FreeSans 200 0 0 0 X
port 7 nsew
flabel pwell s 68 31 102 65 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 68 575 102 609 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 68 31 102 65 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 68 575 102 609 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 38 48 38 48 4 buf_16
<< properties >>
string FIXED_BBOX 38 48 2062 592
string path 0.190 2.960 10.310 2.960 
<< end >>
