magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< pwell >>
rect -26 -26 690 6026
<< nmos >>
rect 132 0 532 6000
<< ndiff >>
rect 0 5969 132 6000
rect 0 5935 13 5969
rect 47 5935 85 5969
rect 119 5935 132 5969
rect 0 5897 132 5935
rect 0 5863 13 5897
rect 47 5863 85 5897
rect 119 5863 132 5897
rect 0 5825 132 5863
rect 0 5791 13 5825
rect 47 5791 85 5825
rect 119 5791 132 5825
rect 0 5753 132 5791
rect 0 5719 13 5753
rect 47 5719 85 5753
rect 119 5719 132 5753
rect 0 5681 132 5719
rect 0 5647 13 5681
rect 47 5647 85 5681
rect 119 5647 132 5681
rect 0 5609 132 5647
rect 0 5575 13 5609
rect 47 5575 85 5609
rect 119 5575 132 5609
rect 0 5537 132 5575
rect 0 5503 13 5537
rect 47 5503 85 5537
rect 119 5503 132 5537
rect 0 5465 132 5503
rect 0 5431 13 5465
rect 47 5431 85 5465
rect 119 5431 132 5465
rect 0 5393 132 5431
rect 0 5359 13 5393
rect 47 5359 85 5393
rect 119 5359 132 5393
rect 0 5321 132 5359
rect 0 5287 13 5321
rect 47 5287 85 5321
rect 119 5287 132 5321
rect 0 5249 132 5287
rect 0 5215 13 5249
rect 47 5215 85 5249
rect 119 5215 132 5249
rect 0 5177 132 5215
rect 0 5143 13 5177
rect 47 5143 85 5177
rect 119 5143 132 5177
rect 0 5105 132 5143
rect 0 5071 13 5105
rect 47 5071 85 5105
rect 119 5071 132 5105
rect 0 5033 132 5071
rect 0 4999 13 5033
rect 47 4999 85 5033
rect 119 4999 132 5033
rect 0 4961 132 4999
rect 0 4927 13 4961
rect 47 4927 85 4961
rect 119 4927 132 4961
rect 0 4889 132 4927
rect 0 4855 13 4889
rect 47 4855 85 4889
rect 119 4855 132 4889
rect 0 4817 132 4855
rect 0 4783 13 4817
rect 47 4783 85 4817
rect 119 4783 132 4817
rect 0 4745 132 4783
rect 0 4711 13 4745
rect 47 4711 85 4745
rect 119 4711 132 4745
rect 0 4673 132 4711
rect 0 4639 13 4673
rect 47 4639 85 4673
rect 119 4639 132 4673
rect 0 4601 132 4639
rect 0 4567 13 4601
rect 47 4567 85 4601
rect 119 4567 132 4601
rect 0 4529 132 4567
rect 0 4495 13 4529
rect 47 4495 85 4529
rect 119 4495 132 4529
rect 0 4457 132 4495
rect 0 4423 13 4457
rect 47 4423 85 4457
rect 119 4423 132 4457
rect 0 4385 132 4423
rect 0 4351 13 4385
rect 47 4351 85 4385
rect 119 4351 132 4385
rect 0 4313 132 4351
rect 0 4279 13 4313
rect 47 4279 85 4313
rect 119 4279 132 4313
rect 0 4241 132 4279
rect 0 4207 13 4241
rect 47 4207 85 4241
rect 119 4207 132 4241
rect 0 4169 132 4207
rect 0 4135 13 4169
rect 47 4135 85 4169
rect 119 4135 132 4169
rect 0 4097 132 4135
rect 0 4063 13 4097
rect 47 4063 85 4097
rect 119 4063 132 4097
rect 0 4025 132 4063
rect 0 3991 13 4025
rect 47 3991 85 4025
rect 119 3991 132 4025
rect 0 3953 132 3991
rect 0 3919 13 3953
rect 47 3919 85 3953
rect 119 3919 132 3953
rect 0 3881 132 3919
rect 0 3847 13 3881
rect 47 3847 85 3881
rect 119 3847 132 3881
rect 0 3809 132 3847
rect 0 3775 13 3809
rect 47 3775 85 3809
rect 119 3775 132 3809
rect 0 3737 132 3775
rect 0 3703 13 3737
rect 47 3703 85 3737
rect 119 3703 132 3737
rect 0 3665 132 3703
rect 0 3631 13 3665
rect 47 3631 85 3665
rect 119 3631 132 3665
rect 0 3593 132 3631
rect 0 3559 13 3593
rect 47 3559 85 3593
rect 119 3559 132 3593
rect 0 3521 132 3559
rect 0 3487 13 3521
rect 47 3487 85 3521
rect 119 3487 132 3521
rect 0 3449 132 3487
rect 0 3415 13 3449
rect 47 3415 85 3449
rect 119 3415 132 3449
rect 0 3377 132 3415
rect 0 3343 13 3377
rect 47 3343 85 3377
rect 119 3343 132 3377
rect 0 3305 132 3343
rect 0 3271 13 3305
rect 47 3271 85 3305
rect 119 3271 132 3305
rect 0 3233 132 3271
rect 0 3199 13 3233
rect 47 3199 85 3233
rect 119 3199 132 3233
rect 0 3161 132 3199
rect 0 3127 13 3161
rect 47 3127 85 3161
rect 119 3127 132 3161
rect 0 3089 132 3127
rect 0 3055 13 3089
rect 47 3055 85 3089
rect 119 3055 132 3089
rect 0 3017 132 3055
rect 0 2983 13 3017
rect 47 2983 85 3017
rect 119 2983 132 3017
rect 0 2945 132 2983
rect 0 2911 13 2945
rect 47 2911 85 2945
rect 119 2911 132 2945
rect 0 2873 132 2911
rect 0 2839 13 2873
rect 47 2839 85 2873
rect 119 2839 132 2873
rect 0 2801 132 2839
rect 0 2767 13 2801
rect 47 2767 85 2801
rect 119 2767 132 2801
rect 0 2729 132 2767
rect 0 2695 13 2729
rect 47 2695 85 2729
rect 119 2695 132 2729
rect 0 2657 132 2695
rect 0 2623 13 2657
rect 47 2623 85 2657
rect 119 2623 132 2657
rect 0 2585 132 2623
rect 0 2551 13 2585
rect 47 2551 85 2585
rect 119 2551 132 2585
rect 0 2513 132 2551
rect 0 2479 13 2513
rect 47 2479 85 2513
rect 119 2479 132 2513
rect 0 2441 132 2479
rect 0 2407 13 2441
rect 47 2407 85 2441
rect 119 2407 132 2441
rect 0 2369 132 2407
rect 0 2335 13 2369
rect 47 2335 85 2369
rect 119 2335 132 2369
rect 0 2297 132 2335
rect 0 2263 13 2297
rect 47 2263 85 2297
rect 119 2263 132 2297
rect 0 2225 132 2263
rect 0 2191 13 2225
rect 47 2191 85 2225
rect 119 2191 132 2225
rect 0 2153 132 2191
rect 0 2119 13 2153
rect 47 2119 85 2153
rect 119 2119 132 2153
rect 0 2081 132 2119
rect 0 2047 13 2081
rect 47 2047 85 2081
rect 119 2047 132 2081
rect 0 2009 132 2047
rect 0 1975 13 2009
rect 47 1975 85 2009
rect 119 1975 132 2009
rect 0 1937 132 1975
rect 0 1903 13 1937
rect 47 1903 85 1937
rect 119 1903 132 1937
rect 0 1865 132 1903
rect 0 1831 13 1865
rect 47 1831 85 1865
rect 119 1831 132 1865
rect 0 1793 132 1831
rect 0 1759 13 1793
rect 47 1759 85 1793
rect 119 1759 132 1793
rect 0 1721 132 1759
rect 0 1687 13 1721
rect 47 1687 85 1721
rect 119 1687 132 1721
rect 0 1649 132 1687
rect 0 1615 13 1649
rect 47 1615 85 1649
rect 119 1615 132 1649
rect 0 1577 132 1615
rect 0 1543 13 1577
rect 47 1543 85 1577
rect 119 1543 132 1577
rect 0 1505 132 1543
rect 0 1471 13 1505
rect 47 1471 85 1505
rect 119 1471 132 1505
rect 0 1433 132 1471
rect 0 1399 13 1433
rect 47 1399 85 1433
rect 119 1399 132 1433
rect 0 1361 132 1399
rect 0 1327 13 1361
rect 47 1327 85 1361
rect 119 1327 132 1361
rect 0 1289 132 1327
rect 0 1255 13 1289
rect 47 1255 85 1289
rect 119 1255 132 1289
rect 0 1217 132 1255
rect 0 1183 13 1217
rect 47 1183 85 1217
rect 119 1183 132 1217
rect 0 1145 132 1183
rect 0 1111 13 1145
rect 47 1111 85 1145
rect 119 1111 132 1145
rect 0 1073 132 1111
rect 0 1039 13 1073
rect 47 1039 85 1073
rect 119 1039 132 1073
rect 0 1001 132 1039
rect 0 967 13 1001
rect 47 967 85 1001
rect 119 967 132 1001
rect 0 929 132 967
rect 0 895 13 929
rect 47 895 85 929
rect 119 895 132 929
rect 0 857 132 895
rect 0 823 13 857
rect 47 823 85 857
rect 119 823 132 857
rect 0 785 132 823
rect 0 751 13 785
rect 47 751 85 785
rect 119 751 132 785
rect 0 713 132 751
rect 0 679 13 713
rect 47 679 85 713
rect 119 679 132 713
rect 0 641 132 679
rect 0 607 13 641
rect 47 607 85 641
rect 119 607 132 641
rect 0 569 132 607
rect 0 535 13 569
rect 47 535 85 569
rect 119 535 132 569
rect 0 497 132 535
rect 0 463 13 497
rect 47 463 85 497
rect 119 463 132 497
rect 0 425 132 463
rect 0 391 13 425
rect 47 391 85 425
rect 119 391 132 425
rect 0 353 132 391
rect 0 319 13 353
rect 47 319 85 353
rect 119 319 132 353
rect 0 281 132 319
rect 0 247 13 281
rect 47 247 85 281
rect 119 247 132 281
rect 0 209 132 247
rect 0 175 13 209
rect 47 175 85 209
rect 119 175 132 209
rect 0 137 132 175
rect 0 103 13 137
rect 47 103 85 137
rect 119 103 132 137
rect 0 65 132 103
rect 0 31 13 65
rect 47 31 85 65
rect 119 31 132 65
rect 0 0 132 31
rect 532 5969 664 6000
rect 532 5935 545 5969
rect 579 5935 617 5969
rect 651 5935 664 5969
rect 532 5897 664 5935
rect 532 5863 545 5897
rect 579 5863 617 5897
rect 651 5863 664 5897
rect 532 5825 664 5863
rect 532 5791 545 5825
rect 579 5791 617 5825
rect 651 5791 664 5825
rect 532 5753 664 5791
rect 532 5719 545 5753
rect 579 5719 617 5753
rect 651 5719 664 5753
rect 532 5681 664 5719
rect 532 5647 545 5681
rect 579 5647 617 5681
rect 651 5647 664 5681
rect 532 5609 664 5647
rect 532 5575 545 5609
rect 579 5575 617 5609
rect 651 5575 664 5609
rect 532 5537 664 5575
rect 532 5503 545 5537
rect 579 5503 617 5537
rect 651 5503 664 5537
rect 532 5465 664 5503
rect 532 5431 545 5465
rect 579 5431 617 5465
rect 651 5431 664 5465
rect 532 5393 664 5431
rect 532 5359 545 5393
rect 579 5359 617 5393
rect 651 5359 664 5393
rect 532 5321 664 5359
rect 532 5287 545 5321
rect 579 5287 617 5321
rect 651 5287 664 5321
rect 532 5249 664 5287
rect 532 5215 545 5249
rect 579 5215 617 5249
rect 651 5215 664 5249
rect 532 5177 664 5215
rect 532 5143 545 5177
rect 579 5143 617 5177
rect 651 5143 664 5177
rect 532 5105 664 5143
rect 532 5071 545 5105
rect 579 5071 617 5105
rect 651 5071 664 5105
rect 532 5033 664 5071
rect 532 4999 545 5033
rect 579 4999 617 5033
rect 651 4999 664 5033
rect 532 4961 664 4999
rect 532 4927 545 4961
rect 579 4927 617 4961
rect 651 4927 664 4961
rect 532 4889 664 4927
rect 532 4855 545 4889
rect 579 4855 617 4889
rect 651 4855 664 4889
rect 532 4817 664 4855
rect 532 4783 545 4817
rect 579 4783 617 4817
rect 651 4783 664 4817
rect 532 4745 664 4783
rect 532 4711 545 4745
rect 579 4711 617 4745
rect 651 4711 664 4745
rect 532 4673 664 4711
rect 532 4639 545 4673
rect 579 4639 617 4673
rect 651 4639 664 4673
rect 532 4601 664 4639
rect 532 4567 545 4601
rect 579 4567 617 4601
rect 651 4567 664 4601
rect 532 4529 664 4567
rect 532 4495 545 4529
rect 579 4495 617 4529
rect 651 4495 664 4529
rect 532 4457 664 4495
rect 532 4423 545 4457
rect 579 4423 617 4457
rect 651 4423 664 4457
rect 532 4385 664 4423
rect 532 4351 545 4385
rect 579 4351 617 4385
rect 651 4351 664 4385
rect 532 4313 664 4351
rect 532 4279 545 4313
rect 579 4279 617 4313
rect 651 4279 664 4313
rect 532 4241 664 4279
rect 532 4207 545 4241
rect 579 4207 617 4241
rect 651 4207 664 4241
rect 532 4169 664 4207
rect 532 4135 545 4169
rect 579 4135 617 4169
rect 651 4135 664 4169
rect 532 4097 664 4135
rect 532 4063 545 4097
rect 579 4063 617 4097
rect 651 4063 664 4097
rect 532 4025 664 4063
rect 532 3991 545 4025
rect 579 3991 617 4025
rect 651 3991 664 4025
rect 532 3953 664 3991
rect 532 3919 545 3953
rect 579 3919 617 3953
rect 651 3919 664 3953
rect 532 3881 664 3919
rect 532 3847 545 3881
rect 579 3847 617 3881
rect 651 3847 664 3881
rect 532 3809 664 3847
rect 532 3775 545 3809
rect 579 3775 617 3809
rect 651 3775 664 3809
rect 532 3737 664 3775
rect 532 3703 545 3737
rect 579 3703 617 3737
rect 651 3703 664 3737
rect 532 3665 664 3703
rect 532 3631 545 3665
rect 579 3631 617 3665
rect 651 3631 664 3665
rect 532 3593 664 3631
rect 532 3559 545 3593
rect 579 3559 617 3593
rect 651 3559 664 3593
rect 532 3521 664 3559
rect 532 3487 545 3521
rect 579 3487 617 3521
rect 651 3487 664 3521
rect 532 3449 664 3487
rect 532 3415 545 3449
rect 579 3415 617 3449
rect 651 3415 664 3449
rect 532 3377 664 3415
rect 532 3343 545 3377
rect 579 3343 617 3377
rect 651 3343 664 3377
rect 532 3305 664 3343
rect 532 3271 545 3305
rect 579 3271 617 3305
rect 651 3271 664 3305
rect 532 3233 664 3271
rect 532 3199 545 3233
rect 579 3199 617 3233
rect 651 3199 664 3233
rect 532 3161 664 3199
rect 532 3127 545 3161
rect 579 3127 617 3161
rect 651 3127 664 3161
rect 532 3089 664 3127
rect 532 3055 545 3089
rect 579 3055 617 3089
rect 651 3055 664 3089
rect 532 3017 664 3055
rect 532 2983 545 3017
rect 579 2983 617 3017
rect 651 2983 664 3017
rect 532 2945 664 2983
rect 532 2911 545 2945
rect 579 2911 617 2945
rect 651 2911 664 2945
rect 532 2873 664 2911
rect 532 2839 545 2873
rect 579 2839 617 2873
rect 651 2839 664 2873
rect 532 2801 664 2839
rect 532 2767 545 2801
rect 579 2767 617 2801
rect 651 2767 664 2801
rect 532 2729 664 2767
rect 532 2695 545 2729
rect 579 2695 617 2729
rect 651 2695 664 2729
rect 532 2657 664 2695
rect 532 2623 545 2657
rect 579 2623 617 2657
rect 651 2623 664 2657
rect 532 2585 664 2623
rect 532 2551 545 2585
rect 579 2551 617 2585
rect 651 2551 664 2585
rect 532 2513 664 2551
rect 532 2479 545 2513
rect 579 2479 617 2513
rect 651 2479 664 2513
rect 532 2441 664 2479
rect 532 2407 545 2441
rect 579 2407 617 2441
rect 651 2407 664 2441
rect 532 2369 664 2407
rect 532 2335 545 2369
rect 579 2335 617 2369
rect 651 2335 664 2369
rect 532 2297 664 2335
rect 532 2263 545 2297
rect 579 2263 617 2297
rect 651 2263 664 2297
rect 532 2225 664 2263
rect 532 2191 545 2225
rect 579 2191 617 2225
rect 651 2191 664 2225
rect 532 2153 664 2191
rect 532 2119 545 2153
rect 579 2119 617 2153
rect 651 2119 664 2153
rect 532 2081 664 2119
rect 532 2047 545 2081
rect 579 2047 617 2081
rect 651 2047 664 2081
rect 532 2009 664 2047
rect 532 1975 545 2009
rect 579 1975 617 2009
rect 651 1975 664 2009
rect 532 1937 664 1975
rect 532 1903 545 1937
rect 579 1903 617 1937
rect 651 1903 664 1937
rect 532 1865 664 1903
rect 532 1831 545 1865
rect 579 1831 617 1865
rect 651 1831 664 1865
rect 532 1793 664 1831
rect 532 1759 545 1793
rect 579 1759 617 1793
rect 651 1759 664 1793
rect 532 1721 664 1759
rect 532 1687 545 1721
rect 579 1687 617 1721
rect 651 1687 664 1721
rect 532 1649 664 1687
rect 532 1615 545 1649
rect 579 1615 617 1649
rect 651 1615 664 1649
rect 532 1577 664 1615
rect 532 1543 545 1577
rect 579 1543 617 1577
rect 651 1543 664 1577
rect 532 1505 664 1543
rect 532 1471 545 1505
rect 579 1471 617 1505
rect 651 1471 664 1505
rect 532 1433 664 1471
rect 532 1399 545 1433
rect 579 1399 617 1433
rect 651 1399 664 1433
rect 532 1361 664 1399
rect 532 1327 545 1361
rect 579 1327 617 1361
rect 651 1327 664 1361
rect 532 1289 664 1327
rect 532 1255 545 1289
rect 579 1255 617 1289
rect 651 1255 664 1289
rect 532 1217 664 1255
rect 532 1183 545 1217
rect 579 1183 617 1217
rect 651 1183 664 1217
rect 532 1145 664 1183
rect 532 1111 545 1145
rect 579 1111 617 1145
rect 651 1111 664 1145
rect 532 1073 664 1111
rect 532 1039 545 1073
rect 579 1039 617 1073
rect 651 1039 664 1073
rect 532 1001 664 1039
rect 532 967 545 1001
rect 579 967 617 1001
rect 651 967 664 1001
rect 532 929 664 967
rect 532 895 545 929
rect 579 895 617 929
rect 651 895 664 929
rect 532 857 664 895
rect 532 823 545 857
rect 579 823 617 857
rect 651 823 664 857
rect 532 785 664 823
rect 532 751 545 785
rect 579 751 617 785
rect 651 751 664 785
rect 532 713 664 751
rect 532 679 545 713
rect 579 679 617 713
rect 651 679 664 713
rect 532 641 664 679
rect 532 607 545 641
rect 579 607 617 641
rect 651 607 664 641
rect 532 569 664 607
rect 532 535 545 569
rect 579 535 617 569
rect 651 535 664 569
rect 532 497 664 535
rect 532 463 545 497
rect 579 463 617 497
rect 651 463 664 497
rect 532 425 664 463
rect 532 391 545 425
rect 579 391 617 425
rect 651 391 664 425
rect 532 353 664 391
rect 532 319 545 353
rect 579 319 617 353
rect 651 319 664 353
rect 532 281 664 319
rect 532 247 545 281
rect 579 247 617 281
rect 651 247 664 281
rect 532 209 664 247
rect 532 175 545 209
rect 579 175 617 209
rect 651 175 664 209
rect 532 137 664 175
rect 532 103 545 137
rect 579 103 617 137
rect 651 103 664 137
rect 532 65 664 103
rect 532 31 545 65
rect 579 31 617 65
rect 651 31 664 65
rect 532 0 664 31
<< ndiffc >>
rect 13 5935 47 5969
rect 85 5935 119 5969
rect 13 5863 47 5897
rect 85 5863 119 5897
rect 13 5791 47 5825
rect 85 5791 119 5825
rect 13 5719 47 5753
rect 85 5719 119 5753
rect 13 5647 47 5681
rect 85 5647 119 5681
rect 13 5575 47 5609
rect 85 5575 119 5609
rect 13 5503 47 5537
rect 85 5503 119 5537
rect 13 5431 47 5465
rect 85 5431 119 5465
rect 13 5359 47 5393
rect 85 5359 119 5393
rect 13 5287 47 5321
rect 85 5287 119 5321
rect 13 5215 47 5249
rect 85 5215 119 5249
rect 13 5143 47 5177
rect 85 5143 119 5177
rect 13 5071 47 5105
rect 85 5071 119 5105
rect 13 4999 47 5033
rect 85 4999 119 5033
rect 13 4927 47 4961
rect 85 4927 119 4961
rect 13 4855 47 4889
rect 85 4855 119 4889
rect 13 4783 47 4817
rect 85 4783 119 4817
rect 13 4711 47 4745
rect 85 4711 119 4745
rect 13 4639 47 4673
rect 85 4639 119 4673
rect 13 4567 47 4601
rect 85 4567 119 4601
rect 13 4495 47 4529
rect 85 4495 119 4529
rect 13 4423 47 4457
rect 85 4423 119 4457
rect 13 4351 47 4385
rect 85 4351 119 4385
rect 13 4279 47 4313
rect 85 4279 119 4313
rect 13 4207 47 4241
rect 85 4207 119 4241
rect 13 4135 47 4169
rect 85 4135 119 4169
rect 13 4063 47 4097
rect 85 4063 119 4097
rect 13 3991 47 4025
rect 85 3991 119 4025
rect 13 3919 47 3953
rect 85 3919 119 3953
rect 13 3847 47 3881
rect 85 3847 119 3881
rect 13 3775 47 3809
rect 85 3775 119 3809
rect 13 3703 47 3737
rect 85 3703 119 3737
rect 13 3631 47 3665
rect 85 3631 119 3665
rect 13 3559 47 3593
rect 85 3559 119 3593
rect 13 3487 47 3521
rect 85 3487 119 3521
rect 13 3415 47 3449
rect 85 3415 119 3449
rect 13 3343 47 3377
rect 85 3343 119 3377
rect 13 3271 47 3305
rect 85 3271 119 3305
rect 13 3199 47 3233
rect 85 3199 119 3233
rect 13 3127 47 3161
rect 85 3127 119 3161
rect 13 3055 47 3089
rect 85 3055 119 3089
rect 13 2983 47 3017
rect 85 2983 119 3017
rect 13 2911 47 2945
rect 85 2911 119 2945
rect 13 2839 47 2873
rect 85 2839 119 2873
rect 13 2767 47 2801
rect 85 2767 119 2801
rect 13 2695 47 2729
rect 85 2695 119 2729
rect 13 2623 47 2657
rect 85 2623 119 2657
rect 13 2551 47 2585
rect 85 2551 119 2585
rect 13 2479 47 2513
rect 85 2479 119 2513
rect 13 2407 47 2441
rect 85 2407 119 2441
rect 13 2335 47 2369
rect 85 2335 119 2369
rect 13 2263 47 2297
rect 85 2263 119 2297
rect 13 2191 47 2225
rect 85 2191 119 2225
rect 13 2119 47 2153
rect 85 2119 119 2153
rect 13 2047 47 2081
rect 85 2047 119 2081
rect 13 1975 47 2009
rect 85 1975 119 2009
rect 13 1903 47 1937
rect 85 1903 119 1937
rect 13 1831 47 1865
rect 85 1831 119 1865
rect 13 1759 47 1793
rect 85 1759 119 1793
rect 13 1687 47 1721
rect 85 1687 119 1721
rect 13 1615 47 1649
rect 85 1615 119 1649
rect 13 1543 47 1577
rect 85 1543 119 1577
rect 13 1471 47 1505
rect 85 1471 119 1505
rect 13 1399 47 1433
rect 85 1399 119 1433
rect 13 1327 47 1361
rect 85 1327 119 1361
rect 13 1255 47 1289
rect 85 1255 119 1289
rect 13 1183 47 1217
rect 85 1183 119 1217
rect 13 1111 47 1145
rect 85 1111 119 1145
rect 13 1039 47 1073
rect 85 1039 119 1073
rect 13 967 47 1001
rect 85 967 119 1001
rect 13 895 47 929
rect 85 895 119 929
rect 13 823 47 857
rect 85 823 119 857
rect 13 751 47 785
rect 85 751 119 785
rect 13 679 47 713
rect 85 679 119 713
rect 13 607 47 641
rect 85 607 119 641
rect 13 535 47 569
rect 85 535 119 569
rect 13 463 47 497
rect 85 463 119 497
rect 13 391 47 425
rect 85 391 119 425
rect 13 319 47 353
rect 85 319 119 353
rect 13 247 47 281
rect 85 247 119 281
rect 13 175 47 209
rect 85 175 119 209
rect 13 103 47 137
rect 85 103 119 137
rect 13 31 47 65
rect 85 31 119 65
rect 545 5935 579 5969
rect 617 5935 651 5969
rect 545 5863 579 5897
rect 617 5863 651 5897
rect 545 5791 579 5825
rect 617 5791 651 5825
rect 545 5719 579 5753
rect 617 5719 651 5753
rect 545 5647 579 5681
rect 617 5647 651 5681
rect 545 5575 579 5609
rect 617 5575 651 5609
rect 545 5503 579 5537
rect 617 5503 651 5537
rect 545 5431 579 5465
rect 617 5431 651 5465
rect 545 5359 579 5393
rect 617 5359 651 5393
rect 545 5287 579 5321
rect 617 5287 651 5321
rect 545 5215 579 5249
rect 617 5215 651 5249
rect 545 5143 579 5177
rect 617 5143 651 5177
rect 545 5071 579 5105
rect 617 5071 651 5105
rect 545 4999 579 5033
rect 617 4999 651 5033
rect 545 4927 579 4961
rect 617 4927 651 4961
rect 545 4855 579 4889
rect 617 4855 651 4889
rect 545 4783 579 4817
rect 617 4783 651 4817
rect 545 4711 579 4745
rect 617 4711 651 4745
rect 545 4639 579 4673
rect 617 4639 651 4673
rect 545 4567 579 4601
rect 617 4567 651 4601
rect 545 4495 579 4529
rect 617 4495 651 4529
rect 545 4423 579 4457
rect 617 4423 651 4457
rect 545 4351 579 4385
rect 617 4351 651 4385
rect 545 4279 579 4313
rect 617 4279 651 4313
rect 545 4207 579 4241
rect 617 4207 651 4241
rect 545 4135 579 4169
rect 617 4135 651 4169
rect 545 4063 579 4097
rect 617 4063 651 4097
rect 545 3991 579 4025
rect 617 3991 651 4025
rect 545 3919 579 3953
rect 617 3919 651 3953
rect 545 3847 579 3881
rect 617 3847 651 3881
rect 545 3775 579 3809
rect 617 3775 651 3809
rect 545 3703 579 3737
rect 617 3703 651 3737
rect 545 3631 579 3665
rect 617 3631 651 3665
rect 545 3559 579 3593
rect 617 3559 651 3593
rect 545 3487 579 3521
rect 617 3487 651 3521
rect 545 3415 579 3449
rect 617 3415 651 3449
rect 545 3343 579 3377
rect 617 3343 651 3377
rect 545 3271 579 3305
rect 617 3271 651 3305
rect 545 3199 579 3233
rect 617 3199 651 3233
rect 545 3127 579 3161
rect 617 3127 651 3161
rect 545 3055 579 3089
rect 617 3055 651 3089
rect 545 2983 579 3017
rect 617 2983 651 3017
rect 545 2911 579 2945
rect 617 2911 651 2945
rect 545 2839 579 2873
rect 617 2839 651 2873
rect 545 2767 579 2801
rect 617 2767 651 2801
rect 545 2695 579 2729
rect 617 2695 651 2729
rect 545 2623 579 2657
rect 617 2623 651 2657
rect 545 2551 579 2585
rect 617 2551 651 2585
rect 545 2479 579 2513
rect 617 2479 651 2513
rect 545 2407 579 2441
rect 617 2407 651 2441
rect 545 2335 579 2369
rect 617 2335 651 2369
rect 545 2263 579 2297
rect 617 2263 651 2297
rect 545 2191 579 2225
rect 617 2191 651 2225
rect 545 2119 579 2153
rect 617 2119 651 2153
rect 545 2047 579 2081
rect 617 2047 651 2081
rect 545 1975 579 2009
rect 617 1975 651 2009
rect 545 1903 579 1937
rect 617 1903 651 1937
rect 545 1831 579 1865
rect 617 1831 651 1865
rect 545 1759 579 1793
rect 617 1759 651 1793
rect 545 1687 579 1721
rect 617 1687 651 1721
rect 545 1615 579 1649
rect 617 1615 651 1649
rect 545 1543 579 1577
rect 617 1543 651 1577
rect 545 1471 579 1505
rect 617 1471 651 1505
rect 545 1399 579 1433
rect 617 1399 651 1433
rect 545 1327 579 1361
rect 617 1327 651 1361
rect 545 1255 579 1289
rect 617 1255 651 1289
rect 545 1183 579 1217
rect 617 1183 651 1217
rect 545 1111 579 1145
rect 617 1111 651 1145
rect 545 1039 579 1073
rect 617 1039 651 1073
rect 545 967 579 1001
rect 617 967 651 1001
rect 545 895 579 929
rect 617 895 651 929
rect 545 823 579 857
rect 617 823 651 857
rect 545 751 579 785
rect 617 751 651 785
rect 545 679 579 713
rect 617 679 651 713
rect 545 607 579 641
rect 617 607 651 641
rect 545 535 579 569
rect 617 535 651 569
rect 545 463 579 497
rect 617 463 651 497
rect 545 391 579 425
rect 617 391 651 425
rect 545 319 579 353
rect 617 319 651 353
rect 545 247 579 281
rect 617 247 651 281
rect 545 175 579 209
rect 617 175 651 209
rect 545 103 579 137
rect 617 103 651 137
rect 545 31 579 65
rect 617 31 651 65
<< poly >>
rect 132 6090 532 6106
rect 132 6056 171 6090
rect 205 6056 243 6090
rect 277 6056 315 6090
rect 349 6056 387 6090
rect 421 6056 459 6090
rect 493 6056 532 6090
rect 132 6000 532 6056
rect 132 -40 532 0
<< polycont >>
rect 171 6056 205 6090
rect 243 6056 277 6090
rect 315 6056 349 6090
rect 387 6056 421 6090
rect 459 6056 493 6090
<< locali >>
rect 155 6056 171 6090
rect 205 6056 243 6090
rect 277 6056 315 6090
rect 349 6056 387 6090
rect 421 6056 459 6090
rect 493 6056 509 6090
rect 13 5969 119 5985
rect 13 15 119 31
rect 545 5969 651 5985
rect 545 15 651 31
<< viali >>
rect 171 6056 205 6090
rect 243 6056 277 6090
rect 315 6056 349 6090
rect 387 6056 421 6090
rect 459 6056 493 6090
rect 13 5935 47 5969
rect 47 5935 85 5969
rect 85 5935 119 5969
rect 13 5897 119 5935
rect 13 5863 47 5897
rect 47 5863 85 5897
rect 85 5863 119 5897
rect 13 5825 119 5863
rect 13 5791 47 5825
rect 47 5791 85 5825
rect 85 5791 119 5825
rect 13 5753 119 5791
rect 13 5719 47 5753
rect 47 5719 85 5753
rect 85 5719 119 5753
rect 13 5681 119 5719
rect 13 5647 47 5681
rect 47 5647 85 5681
rect 85 5647 119 5681
rect 13 5609 119 5647
rect 13 5575 47 5609
rect 47 5575 85 5609
rect 85 5575 119 5609
rect 13 5537 119 5575
rect 13 5503 47 5537
rect 47 5503 85 5537
rect 85 5503 119 5537
rect 13 5465 119 5503
rect 13 5431 47 5465
rect 47 5431 85 5465
rect 85 5431 119 5465
rect 13 5393 119 5431
rect 13 5359 47 5393
rect 47 5359 85 5393
rect 85 5359 119 5393
rect 13 5321 119 5359
rect 13 5287 47 5321
rect 47 5287 85 5321
rect 85 5287 119 5321
rect 13 5249 119 5287
rect 13 5215 47 5249
rect 47 5215 85 5249
rect 85 5215 119 5249
rect 13 5177 119 5215
rect 13 5143 47 5177
rect 47 5143 85 5177
rect 85 5143 119 5177
rect 13 5105 119 5143
rect 13 5071 47 5105
rect 47 5071 85 5105
rect 85 5071 119 5105
rect 13 5033 119 5071
rect 13 4999 47 5033
rect 47 4999 85 5033
rect 85 4999 119 5033
rect 13 4961 119 4999
rect 13 4927 47 4961
rect 47 4927 85 4961
rect 85 4927 119 4961
rect 13 4889 119 4927
rect 13 4855 47 4889
rect 47 4855 85 4889
rect 85 4855 119 4889
rect 13 4817 119 4855
rect 13 4783 47 4817
rect 47 4783 85 4817
rect 85 4783 119 4817
rect 13 4745 119 4783
rect 13 4711 47 4745
rect 47 4711 85 4745
rect 85 4711 119 4745
rect 13 4673 119 4711
rect 13 4639 47 4673
rect 47 4639 85 4673
rect 85 4639 119 4673
rect 13 4601 119 4639
rect 13 4567 47 4601
rect 47 4567 85 4601
rect 85 4567 119 4601
rect 13 4529 119 4567
rect 13 4495 47 4529
rect 47 4495 85 4529
rect 85 4495 119 4529
rect 13 4457 119 4495
rect 13 4423 47 4457
rect 47 4423 85 4457
rect 85 4423 119 4457
rect 13 4385 119 4423
rect 13 4351 47 4385
rect 47 4351 85 4385
rect 85 4351 119 4385
rect 13 4313 119 4351
rect 13 4279 47 4313
rect 47 4279 85 4313
rect 85 4279 119 4313
rect 13 4241 119 4279
rect 13 4207 47 4241
rect 47 4207 85 4241
rect 85 4207 119 4241
rect 13 4169 119 4207
rect 13 4135 47 4169
rect 47 4135 85 4169
rect 85 4135 119 4169
rect 13 4097 119 4135
rect 13 4063 47 4097
rect 47 4063 85 4097
rect 85 4063 119 4097
rect 13 4025 119 4063
rect 13 3991 47 4025
rect 47 3991 85 4025
rect 85 3991 119 4025
rect 13 3953 119 3991
rect 13 3919 47 3953
rect 47 3919 85 3953
rect 85 3919 119 3953
rect 13 3881 119 3919
rect 13 3847 47 3881
rect 47 3847 85 3881
rect 85 3847 119 3881
rect 13 3809 119 3847
rect 13 3775 47 3809
rect 47 3775 85 3809
rect 85 3775 119 3809
rect 13 3737 119 3775
rect 13 3703 47 3737
rect 47 3703 85 3737
rect 85 3703 119 3737
rect 13 3665 119 3703
rect 13 3631 47 3665
rect 47 3631 85 3665
rect 85 3631 119 3665
rect 13 3593 119 3631
rect 13 3559 47 3593
rect 47 3559 85 3593
rect 85 3559 119 3593
rect 13 3521 119 3559
rect 13 3487 47 3521
rect 47 3487 85 3521
rect 85 3487 119 3521
rect 13 3449 119 3487
rect 13 3415 47 3449
rect 47 3415 85 3449
rect 85 3415 119 3449
rect 13 3377 119 3415
rect 13 3343 47 3377
rect 47 3343 85 3377
rect 85 3343 119 3377
rect 13 3305 119 3343
rect 13 3271 47 3305
rect 47 3271 85 3305
rect 85 3271 119 3305
rect 13 3233 119 3271
rect 13 3199 47 3233
rect 47 3199 85 3233
rect 85 3199 119 3233
rect 13 3161 119 3199
rect 13 3127 47 3161
rect 47 3127 85 3161
rect 85 3127 119 3161
rect 13 3089 119 3127
rect 13 3055 47 3089
rect 47 3055 85 3089
rect 85 3055 119 3089
rect 13 3017 119 3055
rect 13 2983 47 3017
rect 47 2983 85 3017
rect 85 2983 119 3017
rect 13 2945 119 2983
rect 13 2911 47 2945
rect 47 2911 85 2945
rect 85 2911 119 2945
rect 13 2873 119 2911
rect 13 2839 47 2873
rect 47 2839 85 2873
rect 85 2839 119 2873
rect 13 2801 119 2839
rect 13 2767 47 2801
rect 47 2767 85 2801
rect 85 2767 119 2801
rect 13 2729 119 2767
rect 13 2695 47 2729
rect 47 2695 85 2729
rect 85 2695 119 2729
rect 13 2657 119 2695
rect 13 2623 47 2657
rect 47 2623 85 2657
rect 85 2623 119 2657
rect 13 2585 119 2623
rect 13 2551 47 2585
rect 47 2551 85 2585
rect 85 2551 119 2585
rect 13 2513 119 2551
rect 13 2479 47 2513
rect 47 2479 85 2513
rect 85 2479 119 2513
rect 13 2441 119 2479
rect 13 2407 47 2441
rect 47 2407 85 2441
rect 85 2407 119 2441
rect 13 2369 119 2407
rect 13 2335 47 2369
rect 47 2335 85 2369
rect 85 2335 119 2369
rect 13 2297 119 2335
rect 13 2263 47 2297
rect 47 2263 85 2297
rect 85 2263 119 2297
rect 13 2225 119 2263
rect 13 2191 47 2225
rect 47 2191 85 2225
rect 85 2191 119 2225
rect 13 2153 119 2191
rect 13 2119 47 2153
rect 47 2119 85 2153
rect 85 2119 119 2153
rect 13 2081 119 2119
rect 13 2047 47 2081
rect 47 2047 85 2081
rect 85 2047 119 2081
rect 13 2009 119 2047
rect 13 1975 47 2009
rect 47 1975 85 2009
rect 85 1975 119 2009
rect 13 1937 119 1975
rect 13 1903 47 1937
rect 47 1903 85 1937
rect 85 1903 119 1937
rect 13 1865 119 1903
rect 13 1831 47 1865
rect 47 1831 85 1865
rect 85 1831 119 1865
rect 13 1793 119 1831
rect 13 1759 47 1793
rect 47 1759 85 1793
rect 85 1759 119 1793
rect 13 1721 119 1759
rect 13 1687 47 1721
rect 47 1687 85 1721
rect 85 1687 119 1721
rect 13 1649 119 1687
rect 13 1615 47 1649
rect 47 1615 85 1649
rect 85 1615 119 1649
rect 13 1577 119 1615
rect 13 1543 47 1577
rect 47 1543 85 1577
rect 85 1543 119 1577
rect 13 1505 119 1543
rect 13 1471 47 1505
rect 47 1471 85 1505
rect 85 1471 119 1505
rect 13 1433 119 1471
rect 13 1399 47 1433
rect 47 1399 85 1433
rect 85 1399 119 1433
rect 13 1361 119 1399
rect 13 1327 47 1361
rect 47 1327 85 1361
rect 85 1327 119 1361
rect 13 1289 119 1327
rect 13 1255 47 1289
rect 47 1255 85 1289
rect 85 1255 119 1289
rect 13 1217 119 1255
rect 13 1183 47 1217
rect 47 1183 85 1217
rect 85 1183 119 1217
rect 13 1145 119 1183
rect 13 1111 47 1145
rect 47 1111 85 1145
rect 85 1111 119 1145
rect 13 1073 119 1111
rect 13 1039 47 1073
rect 47 1039 85 1073
rect 85 1039 119 1073
rect 13 1001 119 1039
rect 13 967 47 1001
rect 47 967 85 1001
rect 85 967 119 1001
rect 13 929 119 967
rect 13 895 47 929
rect 47 895 85 929
rect 85 895 119 929
rect 13 857 119 895
rect 13 823 47 857
rect 47 823 85 857
rect 85 823 119 857
rect 13 785 119 823
rect 13 751 47 785
rect 47 751 85 785
rect 85 751 119 785
rect 13 713 119 751
rect 13 679 47 713
rect 47 679 85 713
rect 85 679 119 713
rect 13 641 119 679
rect 13 607 47 641
rect 47 607 85 641
rect 85 607 119 641
rect 13 569 119 607
rect 13 535 47 569
rect 47 535 85 569
rect 85 535 119 569
rect 13 497 119 535
rect 13 463 47 497
rect 47 463 85 497
rect 85 463 119 497
rect 13 425 119 463
rect 13 391 47 425
rect 47 391 85 425
rect 85 391 119 425
rect 13 353 119 391
rect 13 319 47 353
rect 47 319 85 353
rect 85 319 119 353
rect 13 281 119 319
rect 13 247 47 281
rect 47 247 85 281
rect 85 247 119 281
rect 13 209 119 247
rect 13 175 47 209
rect 47 175 85 209
rect 85 175 119 209
rect 13 137 119 175
rect 13 103 47 137
rect 47 103 85 137
rect 85 103 119 137
rect 13 65 119 103
rect 13 31 47 65
rect 47 31 85 65
rect 85 31 119 65
rect 545 5935 579 5969
rect 579 5935 617 5969
rect 617 5935 651 5969
rect 545 5897 651 5935
rect 545 5863 579 5897
rect 579 5863 617 5897
rect 617 5863 651 5897
rect 545 5825 651 5863
rect 545 5791 579 5825
rect 579 5791 617 5825
rect 617 5791 651 5825
rect 545 5753 651 5791
rect 545 5719 579 5753
rect 579 5719 617 5753
rect 617 5719 651 5753
rect 545 5681 651 5719
rect 545 5647 579 5681
rect 579 5647 617 5681
rect 617 5647 651 5681
rect 545 5609 651 5647
rect 545 5575 579 5609
rect 579 5575 617 5609
rect 617 5575 651 5609
rect 545 5537 651 5575
rect 545 5503 579 5537
rect 579 5503 617 5537
rect 617 5503 651 5537
rect 545 5465 651 5503
rect 545 5431 579 5465
rect 579 5431 617 5465
rect 617 5431 651 5465
rect 545 5393 651 5431
rect 545 5359 579 5393
rect 579 5359 617 5393
rect 617 5359 651 5393
rect 545 5321 651 5359
rect 545 5287 579 5321
rect 579 5287 617 5321
rect 617 5287 651 5321
rect 545 5249 651 5287
rect 545 5215 579 5249
rect 579 5215 617 5249
rect 617 5215 651 5249
rect 545 5177 651 5215
rect 545 5143 579 5177
rect 579 5143 617 5177
rect 617 5143 651 5177
rect 545 5105 651 5143
rect 545 5071 579 5105
rect 579 5071 617 5105
rect 617 5071 651 5105
rect 545 5033 651 5071
rect 545 4999 579 5033
rect 579 4999 617 5033
rect 617 4999 651 5033
rect 545 4961 651 4999
rect 545 4927 579 4961
rect 579 4927 617 4961
rect 617 4927 651 4961
rect 545 4889 651 4927
rect 545 4855 579 4889
rect 579 4855 617 4889
rect 617 4855 651 4889
rect 545 4817 651 4855
rect 545 4783 579 4817
rect 579 4783 617 4817
rect 617 4783 651 4817
rect 545 4745 651 4783
rect 545 4711 579 4745
rect 579 4711 617 4745
rect 617 4711 651 4745
rect 545 4673 651 4711
rect 545 4639 579 4673
rect 579 4639 617 4673
rect 617 4639 651 4673
rect 545 4601 651 4639
rect 545 4567 579 4601
rect 579 4567 617 4601
rect 617 4567 651 4601
rect 545 4529 651 4567
rect 545 4495 579 4529
rect 579 4495 617 4529
rect 617 4495 651 4529
rect 545 4457 651 4495
rect 545 4423 579 4457
rect 579 4423 617 4457
rect 617 4423 651 4457
rect 545 4385 651 4423
rect 545 4351 579 4385
rect 579 4351 617 4385
rect 617 4351 651 4385
rect 545 4313 651 4351
rect 545 4279 579 4313
rect 579 4279 617 4313
rect 617 4279 651 4313
rect 545 4241 651 4279
rect 545 4207 579 4241
rect 579 4207 617 4241
rect 617 4207 651 4241
rect 545 4169 651 4207
rect 545 4135 579 4169
rect 579 4135 617 4169
rect 617 4135 651 4169
rect 545 4097 651 4135
rect 545 4063 579 4097
rect 579 4063 617 4097
rect 617 4063 651 4097
rect 545 4025 651 4063
rect 545 3991 579 4025
rect 579 3991 617 4025
rect 617 3991 651 4025
rect 545 3953 651 3991
rect 545 3919 579 3953
rect 579 3919 617 3953
rect 617 3919 651 3953
rect 545 3881 651 3919
rect 545 3847 579 3881
rect 579 3847 617 3881
rect 617 3847 651 3881
rect 545 3809 651 3847
rect 545 3775 579 3809
rect 579 3775 617 3809
rect 617 3775 651 3809
rect 545 3737 651 3775
rect 545 3703 579 3737
rect 579 3703 617 3737
rect 617 3703 651 3737
rect 545 3665 651 3703
rect 545 3631 579 3665
rect 579 3631 617 3665
rect 617 3631 651 3665
rect 545 3593 651 3631
rect 545 3559 579 3593
rect 579 3559 617 3593
rect 617 3559 651 3593
rect 545 3521 651 3559
rect 545 3487 579 3521
rect 579 3487 617 3521
rect 617 3487 651 3521
rect 545 3449 651 3487
rect 545 3415 579 3449
rect 579 3415 617 3449
rect 617 3415 651 3449
rect 545 3377 651 3415
rect 545 3343 579 3377
rect 579 3343 617 3377
rect 617 3343 651 3377
rect 545 3305 651 3343
rect 545 3271 579 3305
rect 579 3271 617 3305
rect 617 3271 651 3305
rect 545 3233 651 3271
rect 545 3199 579 3233
rect 579 3199 617 3233
rect 617 3199 651 3233
rect 545 3161 651 3199
rect 545 3127 579 3161
rect 579 3127 617 3161
rect 617 3127 651 3161
rect 545 3089 651 3127
rect 545 3055 579 3089
rect 579 3055 617 3089
rect 617 3055 651 3089
rect 545 3017 651 3055
rect 545 2983 579 3017
rect 579 2983 617 3017
rect 617 2983 651 3017
rect 545 2945 651 2983
rect 545 2911 579 2945
rect 579 2911 617 2945
rect 617 2911 651 2945
rect 545 2873 651 2911
rect 545 2839 579 2873
rect 579 2839 617 2873
rect 617 2839 651 2873
rect 545 2801 651 2839
rect 545 2767 579 2801
rect 579 2767 617 2801
rect 617 2767 651 2801
rect 545 2729 651 2767
rect 545 2695 579 2729
rect 579 2695 617 2729
rect 617 2695 651 2729
rect 545 2657 651 2695
rect 545 2623 579 2657
rect 579 2623 617 2657
rect 617 2623 651 2657
rect 545 2585 651 2623
rect 545 2551 579 2585
rect 579 2551 617 2585
rect 617 2551 651 2585
rect 545 2513 651 2551
rect 545 2479 579 2513
rect 579 2479 617 2513
rect 617 2479 651 2513
rect 545 2441 651 2479
rect 545 2407 579 2441
rect 579 2407 617 2441
rect 617 2407 651 2441
rect 545 2369 651 2407
rect 545 2335 579 2369
rect 579 2335 617 2369
rect 617 2335 651 2369
rect 545 2297 651 2335
rect 545 2263 579 2297
rect 579 2263 617 2297
rect 617 2263 651 2297
rect 545 2225 651 2263
rect 545 2191 579 2225
rect 579 2191 617 2225
rect 617 2191 651 2225
rect 545 2153 651 2191
rect 545 2119 579 2153
rect 579 2119 617 2153
rect 617 2119 651 2153
rect 545 2081 651 2119
rect 545 2047 579 2081
rect 579 2047 617 2081
rect 617 2047 651 2081
rect 545 2009 651 2047
rect 545 1975 579 2009
rect 579 1975 617 2009
rect 617 1975 651 2009
rect 545 1937 651 1975
rect 545 1903 579 1937
rect 579 1903 617 1937
rect 617 1903 651 1937
rect 545 1865 651 1903
rect 545 1831 579 1865
rect 579 1831 617 1865
rect 617 1831 651 1865
rect 545 1793 651 1831
rect 545 1759 579 1793
rect 579 1759 617 1793
rect 617 1759 651 1793
rect 545 1721 651 1759
rect 545 1687 579 1721
rect 579 1687 617 1721
rect 617 1687 651 1721
rect 545 1649 651 1687
rect 545 1615 579 1649
rect 579 1615 617 1649
rect 617 1615 651 1649
rect 545 1577 651 1615
rect 545 1543 579 1577
rect 579 1543 617 1577
rect 617 1543 651 1577
rect 545 1505 651 1543
rect 545 1471 579 1505
rect 579 1471 617 1505
rect 617 1471 651 1505
rect 545 1433 651 1471
rect 545 1399 579 1433
rect 579 1399 617 1433
rect 617 1399 651 1433
rect 545 1361 651 1399
rect 545 1327 579 1361
rect 579 1327 617 1361
rect 617 1327 651 1361
rect 545 1289 651 1327
rect 545 1255 579 1289
rect 579 1255 617 1289
rect 617 1255 651 1289
rect 545 1217 651 1255
rect 545 1183 579 1217
rect 579 1183 617 1217
rect 617 1183 651 1217
rect 545 1145 651 1183
rect 545 1111 579 1145
rect 579 1111 617 1145
rect 617 1111 651 1145
rect 545 1073 651 1111
rect 545 1039 579 1073
rect 579 1039 617 1073
rect 617 1039 651 1073
rect 545 1001 651 1039
rect 545 967 579 1001
rect 579 967 617 1001
rect 617 967 651 1001
rect 545 929 651 967
rect 545 895 579 929
rect 579 895 617 929
rect 617 895 651 929
rect 545 857 651 895
rect 545 823 579 857
rect 579 823 617 857
rect 617 823 651 857
rect 545 785 651 823
rect 545 751 579 785
rect 579 751 617 785
rect 617 751 651 785
rect 545 713 651 751
rect 545 679 579 713
rect 579 679 617 713
rect 617 679 651 713
rect 545 641 651 679
rect 545 607 579 641
rect 579 607 617 641
rect 617 607 651 641
rect 545 569 651 607
rect 545 535 579 569
rect 579 535 617 569
rect 617 535 651 569
rect 545 497 651 535
rect 545 463 579 497
rect 579 463 617 497
rect 617 463 651 497
rect 545 425 651 463
rect 545 391 579 425
rect 579 391 617 425
rect 617 391 651 425
rect 545 353 651 391
rect 545 319 579 353
rect 579 319 617 353
rect 617 319 651 353
rect 545 281 651 319
rect 545 247 579 281
rect 579 247 617 281
rect 617 247 651 281
rect 545 209 651 247
rect 545 175 579 209
rect 579 175 617 209
rect 617 175 651 209
rect 545 137 651 175
rect 545 103 579 137
rect 579 103 617 137
rect 617 103 651 137
rect 545 65 651 103
rect 545 31 579 65
rect 579 31 617 65
rect 617 31 651 65
<< metal1 >>
rect 159 6090 505 6096
rect 159 6056 171 6090
rect 205 6056 243 6090
rect 277 6056 315 6090
rect 349 6056 387 6090
rect 421 6056 459 6090
rect 493 6056 505 6090
rect 159 6050 505 6056
rect 7 5969 125 5981
rect 7 31 13 5969
rect 119 31 125 5969
rect 7 19 125 31
rect 539 5969 657 5981
rect 539 31 545 5969
rect 651 31 657 5969
rect 539 19 657 31
<< end >>
