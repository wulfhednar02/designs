magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< xpolycontact >>
rect 92 568 162 1004
rect 92 40 162 476
<< ppolyres >>
rect 92 476 162 568
<< viali >>
rect 110 951 144 985
rect 110 879 144 913
rect 110 807 144 841
rect 110 735 144 769
rect 110 663 144 697
rect 110 591 144 625
rect 110 420 144 454
rect 110 348 144 382
rect 110 276 144 310
rect 110 204 144 238
rect 110 132 144 166
rect 110 60 144 94
<< metal1 >>
rect 102 985 152 998
rect 102 951 110 985
rect 144 951 152 985
rect 102 913 152 951
rect 102 879 110 913
rect 144 879 152 913
rect 102 841 152 879
rect 102 807 110 841
rect 144 807 152 841
rect 102 769 152 807
rect 102 735 110 769
rect 144 735 152 769
rect 102 697 152 735
rect 102 663 110 697
rect 144 663 152 697
rect 102 625 152 663
rect 102 591 110 625
rect 144 591 152 625
rect 102 577 152 591
rect 102 454 152 467
rect 102 420 110 454
rect 144 420 152 454
rect 102 382 152 420
rect 102 348 110 382
rect 144 348 152 382
rect 102 310 152 348
rect 102 276 110 310
rect 144 276 152 310
rect 102 238 152 276
rect 102 204 110 238
rect 144 204 152 238
rect 102 166 152 204
rect 102 132 110 166
rect 144 132 152 166
rect 102 94 152 132
rect 102 60 110 94
rect 144 60 152 94
rect 102 46 152 60
<< end >>
