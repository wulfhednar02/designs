magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< error_s >>
rect -4021 838 2115 881
rect -3953 149 -3715 171
<< viali >>
rect -3930 2151 4024 2329
rect -3922 -105 -3888 -71
rect -3850 -105 -3816 -71
<< metal1 >>
rect -3946 2286 -3939 2338
rect -3887 2329 -3867 2338
rect -3815 2329 -3795 2338
rect -3743 2329 -3723 2338
rect -3671 2329 -3651 2338
rect -3599 2329 -3579 2338
rect -3527 2329 -3507 2338
rect -3455 2329 -3435 2338
rect -3383 2329 -3363 2338
rect -3311 2329 -3291 2338
rect -3239 2329 -3219 2338
rect -3167 2329 -3147 2338
rect -3095 2329 -3075 2338
rect -3023 2329 -3003 2338
rect -2951 2329 -2931 2338
rect -2879 2329 -2859 2338
rect -2807 2329 -2787 2338
rect -2735 2329 -2715 2338
rect -2663 2329 -2643 2338
rect -2591 2329 -2571 2338
rect -2519 2329 -2499 2338
rect -2447 2329 -2427 2338
rect -2375 2329 -2355 2338
rect -2303 2329 -2283 2338
rect -2231 2329 -2211 2338
rect -2159 2329 -2139 2338
rect -2087 2329 -2067 2338
rect -2015 2329 -1995 2338
rect -1943 2329 -1923 2338
rect -1871 2329 -1851 2338
rect -1799 2329 -1779 2338
rect -1727 2329 -1707 2338
rect -1655 2329 -1635 2338
rect -1583 2329 -1563 2338
rect -1511 2329 -1491 2338
rect -1439 2329 -1419 2338
rect -1367 2329 -1347 2338
rect -1295 2329 -1275 2338
rect -1223 2329 -1203 2338
rect -1151 2329 -1131 2338
rect -1079 2329 -1059 2338
rect -1007 2329 -987 2338
rect -935 2329 -915 2338
rect -863 2329 -843 2338
rect -791 2329 -771 2338
rect -719 2329 -699 2338
rect -647 2329 -627 2338
rect -575 2329 -555 2338
rect -503 2329 -483 2338
rect -431 2329 -411 2338
rect -359 2329 -339 2338
rect -287 2329 -267 2338
rect -215 2329 -195 2338
rect -143 2329 -123 2338
rect -71 2329 -51 2338
rect 1 2329 21 2338
rect 73 2329 93 2338
rect 145 2329 165 2338
rect 217 2329 237 2338
rect 289 2329 309 2338
rect 361 2329 381 2338
rect 433 2329 453 2338
rect 505 2329 525 2338
rect 577 2329 597 2338
rect 649 2329 669 2338
rect 721 2329 741 2338
rect 793 2329 813 2338
rect 865 2329 885 2338
rect 937 2329 957 2338
rect 1009 2329 1029 2338
rect 1081 2329 1101 2338
rect 1153 2329 1173 2338
rect 1225 2329 1245 2338
rect 1297 2329 1317 2338
rect 1369 2329 1389 2338
rect 1441 2329 1461 2338
rect 1513 2329 1533 2338
rect 1585 2329 1605 2338
rect 1657 2329 1677 2338
rect 1729 2329 1749 2338
rect 1801 2329 1821 2338
rect 1873 2329 1893 2338
rect 1945 2329 1965 2338
rect 2017 2329 2037 2338
rect 2089 2329 2109 2338
rect 2161 2329 2181 2338
rect 2233 2329 2253 2338
rect 2305 2329 2325 2338
rect 2377 2329 2397 2338
rect 2449 2329 2469 2338
rect 2521 2329 2541 2338
rect 2593 2329 2613 2338
rect 2665 2329 2685 2338
rect 2737 2329 2757 2338
rect 2809 2329 2829 2338
rect 2881 2329 2901 2338
rect 2953 2329 2973 2338
rect 3025 2329 3045 2338
rect 3097 2329 3117 2338
rect 3169 2329 3189 2338
rect 3241 2329 3261 2338
rect 3313 2329 3333 2338
rect 3385 2329 3405 2338
rect 3457 2329 3477 2338
rect 3529 2329 3549 2338
rect 3601 2329 3621 2338
rect 3673 2329 3693 2338
rect 3745 2329 3765 2338
rect 3817 2329 3837 2338
rect 3889 2329 3909 2338
rect 3961 2329 3981 2338
rect 4033 2286 4040 2338
rect -3946 2266 -3930 2286
rect 4024 2266 4040 2286
rect -3946 2214 -3939 2266
rect 4033 2214 4040 2266
rect -3946 2194 -3930 2214
rect 4024 2194 4040 2214
rect -3946 2151 -3939 2194
rect 4033 2151 4040 2194
rect -3942 2142 -3939 2151
rect -3887 2142 -3867 2151
rect -3815 2142 -3795 2151
rect -3743 2142 -3723 2151
rect -3671 2142 -3651 2151
rect -3599 2142 -3579 2151
rect -3527 2142 -3507 2151
rect -3455 2142 -3435 2151
rect -3383 2142 -3363 2151
rect -3311 2142 -3291 2151
rect -3239 2142 -3219 2151
rect -3167 2142 -3147 2151
rect -3095 2142 -3075 2151
rect -3023 2142 -3003 2151
rect -2951 2142 -2931 2151
rect -2879 2142 -2859 2151
rect -2807 2142 -2787 2151
rect -2735 2142 -2715 2151
rect -2663 2142 -2643 2151
rect -2591 2142 -2571 2151
rect -2519 2142 -2499 2151
rect -2447 2142 -2427 2151
rect -2375 2142 -2355 2151
rect -2303 2142 -2283 2151
rect -2231 2142 -2211 2151
rect -2159 2142 -2139 2151
rect -2087 2142 -2067 2151
rect -2015 2142 -1995 2151
rect -1943 2142 -1923 2151
rect -1871 2142 -1851 2151
rect -1799 2142 -1779 2151
rect -1727 2142 -1707 2151
rect -1655 2142 -1635 2151
rect -1583 2142 -1563 2151
rect -1511 2142 -1491 2151
rect -1439 2142 -1419 2151
rect -1367 2142 -1347 2151
rect -1295 2142 -1275 2151
rect -1223 2142 -1203 2151
rect -1151 2142 -1131 2151
rect -1079 2142 -1059 2151
rect -1007 2142 -987 2151
rect -935 2142 -915 2151
rect -863 2142 -843 2151
rect -791 2142 -771 2151
rect -719 2142 -699 2151
rect -647 2142 -627 2151
rect -575 2142 -555 2151
rect -503 2142 -483 2151
rect -431 2142 -411 2151
rect -359 2142 -339 2151
rect -287 2142 -267 2151
rect -215 2142 -195 2151
rect -143 2142 -123 2151
rect -71 2142 -51 2151
rect 1 2142 21 2151
rect 73 2142 93 2151
rect 145 2142 165 2151
rect 217 2142 237 2151
rect 289 2142 309 2151
rect 361 2142 381 2151
rect 433 2142 453 2151
rect 505 2142 525 2151
rect 577 2142 597 2151
rect 649 2142 669 2151
rect 721 2142 741 2151
rect 793 2142 813 2151
rect 865 2142 885 2151
rect 937 2142 957 2151
rect 1009 2142 1029 2151
rect 1081 2142 1101 2151
rect 1153 2142 1173 2151
rect 1225 2142 1245 2151
rect 1297 2142 1317 2151
rect 1369 2142 1389 2151
rect 1441 2142 1461 2151
rect 1513 2142 1533 2151
rect 1585 2142 1605 2151
rect 1657 2142 1677 2151
rect 1729 2142 1749 2151
rect 1801 2142 1821 2151
rect 1873 2142 1893 2151
rect 1945 2142 1965 2151
rect 2017 2142 2037 2151
rect 2089 2142 2109 2151
rect 2161 2142 2181 2151
rect 2233 2142 2253 2151
rect 2305 2142 2325 2151
rect 2377 2142 2397 2151
rect 2449 2142 2469 2151
rect 2521 2142 2541 2151
rect 2593 2142 2613 2151
rect 2665 2142 2685 2151
rect 2737 2142 2757 2151
rect 2809 2142 2829 2151
rect 2881 2142 2901 2151
rect 2953 2142 2973 2151
rect 3025 2142 3045 2151
rect 3097 2142 3117 2151
rect 3169 2142 3189 2151
rect 3241 2142 3261 2151
rect 3313 2142 3333 2151
rect 3385 2142 3405 2151
rect 3457 2142 3477 2151
rect 3529 2142 3549 2151
rect 3601 2142 3621 2151
rect 3673 2142 3693 2151
rect 3745 2142 3765 2151
rect 3817 2142 3837 2151
rect 3889 2142 3909 2151
rect 3961 2142 3981 2151
rect 4033 2142 4036 2151
rect -3942 2100 4036 2142
rect -4118 308 -4003 1892
rect -3942 688 4036 1096
rect -4110 -31 -3974 105
rect -3938 64 -3800 274
rect -3938 4 -3800 10
rect -3938 -48 -3932 4
rect -3880 -48 -3858 4
rect -3806 -48 -3800 4
rect -3938 -70 -3800 -48
rect -3938 -122 -3932 -70
rect -3880 -122 -3858 -70
rect -3806 -122 -3800 -70
rect -3938 -128 -3800 -122
<< via1 >>
rect -3939 2329 -3887 2338
rect -3867 2329 -3815 2338
rect -3795 2329 -3743 2338
rect -3723 2329 -3671 2338
rect -3651 2329 -3599 2338
rect -3579 2329 -3527 2338
rect -3507 2329 -3455 2338
rect -3435 2329 -3383 2338
rect -3363 2329 -3311 2338
rect -3291 2329 -3239 2338
rect -3219 2329 -3167 2338
rect -3147 2329 -3095 2338
rect -3075 2329 -3023 2338
rect -3003 2329 -2951 2338
rect -2931 2329 -2879 2338
rect -2859 2329 -2807 2338
rect -2787 2329 -2735 2338
rect -2715 2329 -2663 2338
rect -2643 2329 -2591 2338
rect -2571 2329 -2519 2338
rect -2499 2329 -2447 2338
rect -2427 2329 -2375 2338
rect -2355 2329 -2303 2338
rect -2283 2329 -2231 2338
rect -2211 2329 -2159 2338
rect -2139 2329 -2087 2338
rect -2067 2329 -2015 2338
rect -1995 2329 -1943 2338
rect -1923 2329 -1871 2338
rect -1851 2329 -1799 2338
rect -1779 2329 -1727 2338
rect -1707 2329 -1655 2338
rect -1635 2329 -1583 2338
rect -1563 2329 -1511 2338
rect -1491 2329 -1439 2338
rect -1419 2329 -1367 2338
rect -1347 2329 -1295 2338
rect -1275 2329 -1223 2338
rect -1203 2329 -1151 2338
rect -1131 2329 -1079 2338
rect -1059 2329 -1007 2338
rect -987 2329 -935 2338
rect -915 2329 -863 2338
rect -843 2329 -791 2338
rect -771 2329 -719 2338
rect -699 2329 -647 2338
rect -627 2329 -575 2338
rect -555 2329 -503 2338
rect -483 2329 -431 2338
rect -411 2329 -359 2338
rect -339 2329 -287 2338
rect -267 2329 -215 2338
rect -195 2329 -143 2338
rect -123 2329 -71 2338
rect -51 2329 1 2338
rect 21 2329 73 2338
rect 93 2329 145 2338
rect 165 2329 217 2338
rect 237 2329 289 2338
rect 309 2329 361 2338
rect 381 2329 433 2338
rect 453 2329 505 2338
rect 525 2329 577 2338
rect 597 2329 649 2338
rect 669 2329 721 2338
rect 741 2329 793 2338
rect 813 2329 865 2338
rect 885 2329 937 2338
rect 957 2329 1009 2338
rect 1029 2329 1081 2338
rect 1101 2329 1153 2338
rect 1173 2329 1225 2338
rect 1245 2329 1297 2338
rect 1317 2329 1369 2338
rect 1389 2329 1441 2338
rect 1461 2329 1513 2338
rect 1533 2329 1585 2338
rect 1605 2329 1657 2338
rect 1677 2329 1729 2338
rect 1749 2329 1801 2338
rect 1821 2329 1873 2338
rect 1893 2329 1945 2338
rect 1965 2329 2017 2338
rect 2037 2329 2089 2338
rect 2109 2329 2161 2338
rect 2181 2329 2233 2338
rect 2253 2329 2305 2338
rect 2325 2329 2377 2338
rect 2397 2329 2449 2338
rect 2469 2329 2521 2338
rect 2541 2329 2593 2338
rect 2613 2329 2665 2338
rect 2685 2329 2737 2338
rect 2757 2329 2809 2338
rect 2829 2329 2881 2338
rect 2901 2329 2953 2338
rect 2973 2329 3025 2338
rect 3045 2329 3097 2338
rect 3117 2329 3169 2338
rect 3189 2329 3241 2338
rect 3261 2329 3313 2338
rect 3333 2329 3385 2338
rect 3405 2329 3457 2338
rect 3477 2329 3529 2338
rect 3549 2329 3601 2338
rect 3621 2329 3673 2338
rect 3693 2329 3745 2338
rect 3765 2329 3817 2338
rect 3837 2329 3889 2338
rect 3909 2329 3961 2338
rect 3981 2329 4033 2338
rect -3939 2286 -3930 2329
rect -3930 2286 -3887 2329
rect -3867 2286 -3815 2329
rect -3795 2286 -3743 2329
rect -3723 2286 -3671 2329
rect -3651 2286 -3599 2329
rect -3579 2286 -3527 2329
rect -3507 2286 -3455 2329
rect -3435 2286 -3383 2329
rect -3363 2286 -3311 2329
rect -3291 2286 -3239 2329
rect -3219 2286 -3167 2329
rect -3147 2286 -3095 2329
rect -3075 2286 -3023 2329
rect -3003 2286 -2951 2329
rect -2931 2286 -2879 2329
rect -2859 2286 -2807 2329
rect -2787 2286 -2735 2329
rect -2715 2286 -2663 2329
rect -2643 2286 -2591 2329
rect -2571 2286 -2519 2329
rect -2499 2286 -2447 2329
rect -2427 2286 -2375 2329
rect -2355 2286 -2303 2329
rect -2283 2286 -2231 2329
rect -2211 2286 -2159 2329
rect -2139 2286 -2087 2329
rect -2067 2286 -2015 2329
rect -1995 2286 -1943 2329
rect -1923 2286 -1871 2329
rect -1851 2286 -1799 2329
rect -1779 2286 -1727 2329
rect -1707 2286 -1655 2329
rect -1635 2286 -1583 2329
rect -1563 2286 -1511 2329
rect -1491 2286 -1439 2329
rect -1419 2286 -1367 2329
rect -1347 2286 -1295 2329
rect -1275 2286 -1223 2329
rect -1203 2286 -1151 2329
rect -1131 2286 -1079 2329
rect -1059 2286 -1007 2329
rect -987 2286 -935 2329
rect -915 2286 -863 2329
rect -843 2286 -791 2329
rect -771 2286 -719 2329
rect -699 2286 -647 2329
rect -627 2286 -575 2329
rect -555 2286 -503 2329
rect -483 2286 -431 2329
rect -411 2286 -359 2329
rect -339 2286 -287 2329
rect -267 2286 -215 2329
rect -195 2286 -143 2329
rect -123 2286 -71 2329
rect -51 2286 1 2329
rect 21 2286 73 2329
rect 93 2286 145 2329
rect 165 2286 217 2329
rect 237 2286 289 2329
rect 309 2286 361 2329
rect 381 2286 433 2329
rect 453 2286 505 2329
rect 525 2286 577 2329
rect 597 2286 649 2329
rect 669 2286 721 2329
rect 741 2286 793 2329
rect 813 2286 865 2329
rect 885 2286 937 2329
rect 957 2286 1009 2329
rect 1029 2286 1081 2329
rect 1101 2286 1153 2329
rect 1173 2286 1225 2329
rect 1245 2286 1297 2329
rect 1317 2286 1369 2329
rect 1389 2286 1441 2329
rect 1461 2286 1513 2329
rect 1533 2286 1585 2329
rect 1605 2286 1657 2329
rect 1677 2286 1729 2329
rect 1749 2286 1801 2329
rect 1821 2286 1873 2329
rect 1893 2286 1945 2329
rect 1965 2286 2017 2329
rect 2037 2286 2089 2329
rect 2109 2286 2161 2329
rect 2181 2286 2233 2329
rect 2253 2286 2305 2329
rect 2325 2286 2377 2329
rect 2397 2286 2449 2329
rect 2469 2286 2521 2329
rect 2541 2286 2593 2329
rect 2613 2286 2665 2329
rect 2685 2286 2737 2329
rect 2757 2286 2809 2329
rect 2829 2286 2881 2329
rect 2901 2286 2953 2329
rect 2973 2286 3025 2329
rect 3045 2286 3097 2329
rect 3117 2286 3169 2329
rect 3189 2286 3241 2329
rect 3261 2286 3313 2329
rect 3333 2286 3385 2329
rect 3405 2286 3457 2329
rect 3477 2286 3529 2329
rect 3549 2286 3601 2329
rect 3621 2286 3673 2329
rect 3693 2286 3745 2329
rect 3765 2286 3817 2329
rect 3837 2286 3889 2329
rect 3909 2286 3961 2329
rect 3981 2286 4024 2329
rect 4024 2286 4033 2329
rect -3939 2214 -3930 2266
rect -3930 2214 -3887 2266
rect -3867 2214 -3815 2266
rect -3795 2214 -3743 2266
rect -3723 2214 -3671 2266
rect -3651 2214 -3599 2266
rect -3579 2214 -3527 2266
rect -3507 2214 -3455 2266
rect -3435 2214 -3383 2266
rect -3363 2214 -3311 2266
rect -3291 2214 -3239 2266
rect -3219 2214 -3167 2266
rect -3147 2214 -3095 2266
rect -3075 2214 -3023 2266
rect -3003 2214 -2951 2266
rect -2931 2214 -2879 2266
rect -2859 2214 -2807 2266
rect -2787 2214 -2735 2266
rect -2715 2214 -2663 2266
rect -2643 2214 -2591 2266
rect -2571 2214 -2519 2266
rect -2499 2214 -2447 2266
rect -2427 2214 -2375 2266
rect -2355 2214 -2303 2266
rect -2283 2214 -2231 2266
rect -2211 2214 -2159 2266
rect -2139 2214 -2087 2266
rect -2067 2214 -2015 2266
rect -1995 2214 -1943 2266
rect -1923 2214 -1871 2266
rect -1851 2214 -1799 2266
rect -1779 2214 -1727 2266
rect -1707 2214 -1655 2266
rect -1635 2214 -1583 2266
rect -1563 2214 -1511 2266
rect -1491 2214 -1439 2266
rect -1419 2214 -1367 2266
rect -1347 2214 -1295 2266
rect -1275 2214 -1223 2266
rect -1203 2214 -1151 2266
rect -1131 2214 -1079 2266
rect -1059 2214 -1007 2266
rect -987 2214 -935 2266
rect -915 2214 -863 2266
rect -843 2214 -791 2266
rect -771 2214 -719 2266
rect -699 2214 -647 2266
rect -627 2214 -575 2266
rect -555 2214 -503 2266
rect -483 2214 -431 2266
rect -411 2214 -359 2266
rect -339 2214 -287 2266
rect -267 2214 -215 2266
rect -195 2214 -143 2266
rect -123 2214 -71 2266
rect -51 2214 1 2266
rect 21 2214 73 2266
rect 93 2214 145 2266
rect 165 2214 217 2266
rect 237 2214 289 2266
rect 309 2214 361 2266
rect 381 2214 433 2266
rect 453 2214 505 2266
rect 525 2214 577 2266
rect 597 2214 649 2266
rect 669 2214 721 2266
rect 741 2214 793 2266
rect 813 2214 865 2266
rect 885 2214 937 2266
rect 957 2214 1009 2266
rect 1029 2214 1081 2266
rect 1101 2214 1153 2266
rect 1173 2214 1225 2266
rect 1245 2214 1297 2266
rect 1317 2214 1369 2266
rect 1389 2214 1441 2266
rect 1461 2214 1513 2266
rect 1533 2214 1585 2266
rect 1605 2214 1657 2266
rect 1677 2214 1729 2266
rect 1749 2214 1801 2266
rect 1821 2214 1873 2266
rect 1893 2214 1945 2266
rect 1965 2214 2017 2266
rect 2037 2214 2089 2266
rect 2109 2214 2161 2266
rect 2181 2214 2233 2266
rect 2253 2214 2305 2266
rect 2325 2214 2377 2266
rect 2397 2214 2449 2266
rect 2469 2214 2521 2266
rect 2541 2214 2593 2266
rect 2613 2214 2665 2266
rect 2685 2214 2737 2266
rect 2757 2214 2809 2266
rect 2829 2214 2881 2266
rect 2901 2214 2953 2266
rect 2973 2214 3025 2266
rect 3045 2214 3097 2266
rect 3117 2214 3169 2266
rect 3189 2214 3241 2266
rect 3261 2214 3313 2266
rect 3333 2214 3385 2266
rect 3405 2214 3457 2266
rect 3477 2214 3529 2266
rect 3549 2214 3601 2266
rect 3621 2214 3673 2266
rect 3693 2214 3745 2266
rect 3765 2214 3817 2266
rect 3837 2214 3889 2266
rect 3909 2214 3961 2266
rect 3981 2214 4024 2266
rect 4024 2214 4033 2266
rect -3939 2151 -3930 2194
rect -3930 2151 -3887 2194
rect -3867 2151 -3815 2194
rect -3795 2151 -3743 2194
rect -3723 2151 -3671 2194
rect -3651 2151 -3599 2194
rect -3579 2151 -3527 2194
rect -3507 2151 -3455 2194
rect -3435 2151 -3383 2194
rect -3363 2151 -3311 2194
rect -3291 2151 -3239 2194
rect -3219 2151 -3167 2194
rect -3147 2151 -3095 2194
rect -3075 2151 -3023 2194
rect -3003 2151 -2951 2194
rect -2931 2151 -2879 2194
rect -2859 2151 -2807 2194
rect -2787 2151 -2735 2194
rect -2715 2151 -2663 2194
rect -2643 2151 -2591 2194
rect -2571 2151 -2519 2194
rect -2499 2151 -2447 2194
rect -2427 2151 -2375 2194
rect -2355 2151 -2303 2194
rect -2283 2151 -2231 2194
rect -2211 2151 -2159 2194
rect -2139 2151 -2087 2194
rect -2067 2151 -2015 2194
rect -1995 2151 -1943 2194
rect -1923 2151 -1871 2194
rect -1851 2151 -1799 2194
rect -1779 2151 -1727 2194
rect -1707 2151 -1655 2194
rect -1635 2151 -1583 2194
rect -1563 2151 -1511 2194
rect -1491 2151 -1439 2194
rect -1419 2151 -1367 2194
rect -1347 2151 -1295 2194
rect -1275 2151 -1223 2194
rect -1203 2151 -1151 2194
rect -1131 2151 -1079 2194
rect -1059 2151 -1007 2194
rect -987 2151 -935 2194
rect -915 2151 -863 2194
rect -843 2151 -791 2194
rect -771 2151 -719 2194
rect -699 2151 -647 2194
rect -627 2151 -575 2194
rect -555 2151 -503 2194
rect -483 2151 -431 2194
rect -411 2151 -359 2194
rect -339 2151 -287 2194
rect -267 2151 -215 2194
rect -195 2151 -143 2194
rect -123 2151 -71 2194
rect -51 2151 1 2194
rect 21 2151 73 2194
rect 93 2151 145 2194
rect 165 2151 217 2194
rect 237 2151 289 2194
rect 309 2151 361 2194
rect 381 2151 433 2194
rect 453 2151 505 2194
rect 525 2151 577 2194
rect 597 2151 649 2194
rect 669 2151 721 2194
rect 741 2151 793 2194
rect 813 2151 865 2194
rect 885 2151 937 2194
rect 957 2151 1009 2194
rect 1029 2151 1081 2194
rect 1101 2151 1153 2194
rect 1173 2151 1225 2194
rect 1245 2151 1297 2194
rect 1317 2151 1369 2194
rect 1389 2151 1441 2194
rect 1461 2151 1513 2194
rect 1533 2151 1585 2194
rect 1605 2151 1657 2194
rect 1677 2151 1729 2194
rect 1749 2151 1801 2194
rect 1821 2151 1873 2194
rect 1893 2151 1945 2194
rect 1965 2151 2017 2194
rect 2037 2151 2089 2194
rect 2109 2151 2161 2194
rect 2181 2151 2233 2194
rect 2253 2151 2305 2194
rect 2325 2151 2377 2194
rect 2397 2151 2449 2194
rect 2469 2151 2521 2194
rect 2541 2151 2593 2194
rect 2613 2151 2665 2194
rect 2685 2151 2737 2194
rect 2757 2151 2809 2194
rect 2829 2151 2881 2194
rect 2901 2151 2953 2194
rect 2973 2151 3025 2194
rect 3045 2151 3097 2194
rect 3117 2151 3169 2194
rect 3189 2151 3241 2194
rect 3261 2151 3313 2194
rect 3333 2151 3385 2194
rect 3405 2151 3457 2194
rect 3477 2151 3529 2194
rect 3549 2151 3601 2194
rect 3621 2151 3673 2194
rect 3693 2151 3745 2194
rect 3765 2151 3817 2194
rect 3837 2151 3889 2194
rect 3909 2151 3961 2194
rect 3981 2151 4024 2194
rect 4024 2151 4033 2194
rect -3939 2142 -3887 2151
rect -3867 2142 -3815 2151
rect -3795 2142 -3743 2151
rect -3723 2142 -3671 2151
rect -3651 2142 -3599 2151
rect -3579 2142 -3527 2151
rect -3507 2142 -3455 2151
rect -3435 2142 -3383 2151
rect -3363 2142 -3311 2151
rect -3291 2142 -3239 2151
rect -3219 2142 -3167 2151
rect -3147 2142 -3095 2151
rect -3075 2142 -3023 2151
rect -3003 2142 -2951 2151
rect -2931 2142 -2879 2151
rect -2859 2142 -2807 2151
rect -2787 2142 -2735 2151
rect -2715 2142 -2663 2151
rect -2643 2142 -2591 2151
rect -2571 2142 -2519 2151
rect -2499 2142 -2447 2151
rect -2427 2142 -2375 2151
rect -2355 2142 -2303 2151
rect -2283 2142 -2231 2151
rect -2211 2142 -2159 2151
rect -2139 2142 -2087 2151
rect -2067 2142 -2015 2151
rect -1995 2142 -1943 2151
rect -1923 2142 -1871 2151
rect -1851 2142 -1799 2151
rect -1779 2142 -1727 2151
rect -1707 2142 -1655 2151
rect -1635 2142 -1583 2151
rect -1563 2142 -1511 2151
rect -1491 2142 -1439 2151
rect -1419 2142 -1367 2151
rect -1347 2142 -1295 2151
rect -1275 2142 -1223 2151
rect -1203 2142 -1151 2151
rect -1131 2142 -1079 2151
rect -1059 2142 -1007 2151
rect -987 2142 -935 2151
rect -915 2142 -863 2151
rect -843 2142 -791 2151
rect -771 2142 -719 2151
rect -699 2142 -647 2151
rect -627 2142 -575 2151
rect -555 2142 -503 2151
rect -483 2142 -431 2151
rect -411 2142 -359 2151
rect -339 2142 -287 2151
rect -267 2142 -215 2151
rect -195 2142 -143 2151
rect -123 2142 -71 2151
rect -51 2142 1 2151
rect 21 2142 73 2151
rect 93 2142 145 2151
rect 165 2142 217 2151
rect 237 2142 289 2151
rect 309 2142 361 2151
rect 381 2142 433 2151
rect 453 2142 505 2151
rect 525 2142 577 2151
rect 597 2142 649 2151
rect 669 2142 721 2151
rect 741 2142 793 2151
rect 813 2142 865 2151
rect 885 2142 937 2151
rect 957 2142 1009 2151
rect 1029 2142 1081 2151
rect 1101 2142 1153 2151
rect 1173 2142 1225 2151
rect 1245 2142 1297 2151
rect 1317 2142 1369 2151
rect 1389 2142 1441 2151
rect 1461 2142 1513 2151
rect 1533 2142 1585 2151
rect 1605 2142 1657 2151
rect 1677 2142 1729 2151
rect 1749 2142 1801 2151
rect 1821 2142 1873 2151
rect 1893 2142 1945 2151
rect 1965 2142 2017 2151
rect 2037 2142 2089 2151
rect 2109 2142 2161 2151
rect 2181 2142 2233 2151
rect 2253 2142 2305 2151
rect 2325 2142 2377 2151
rect 2397 2142 2449 2151
rect 2469 2142 2521 2151
rect 2541 2142 2593 2151
rect 2613 2142 2665 2151
rect 2685 2142 2737 2151
rect 2757 2142 2809 2151
rect 2829 2142 2881 2151
rect 2901 2142 2953 2151
rect 2973 2142 3025 2151
rect 3045 2142 3097 2151
rect 3117 2142 3169 2151
rect 3189 2142 3241 2151
rect 3261 2142 3313 2151
rect 3333 2142 3385 2151
rect 3405 2142 3457 2151
rect 3477 2142 3529 2151
rect 3549 2142 3601 2151
rect 3621 2142 3673 2151
rect 3693 2142 3745 2151
rect 3765 2142 3817 2151
rect 3837 2142 3889 2151
rect 3909 2142 3961 2151
rect 3981 2142 4033 2151
rect -3932 -48 -3880 4
rect -3858 -48 -3806 4
rect -3932 -71 -3880 -70
rect -3932 -105 -3922 -71
rect -3922 -105 -3888 -71
rect -3888 -105 -3880 -71
rect -3932 -122 -3880 -105
rect -3858 -71 -3806 -70
rect -3858 -105 -3850 -71
rect -3850 -105 -3816 -71
rect -3816 -105 -3806 -71
rect -3858 -122 -3806 -105
<< metal2 >>
rect -3945 2338 4039 2344
rect -3945 2286 -3939 2338
rect -3887 2286 -3867 2338
rect -3815 2286 -3795 2338
rect -3743 2286 -3723 2338
rect -3671 2286 -3651 2338
rect -3599 2286 -3579 2338
rect -3527 2286 -3507 2338
rect -3455 2286 -3435 2338
rect -3383 2286 -3363 2338
rect -3311 2286 -3291 2338
rect -3239 2286 -3219 2338
rect -3167 2286 -3147 2338
rect -3095 2286 -3075 2338
rect -3023 2286 -3003 2338
rect -2951 2286 -2931 2338
rect -2879 2286 -2859 2338
rect -2807 2286 -2787 2338
rect -2735 2286 -2715 2338
rect -2663 2286 -2643 2338
rect -2591 2286 -2571 2338
rect -2519 2286 -2499 2338
rect -2447 2286 -2427 2338
rect -2375 2286 -2355 2338
rect -2303 2286 -2283 2338
rect -2231 2286 -2211 2338
rect -2159 2286 -2139 2338
rect -2087 2286 -2067 2338
rect -2015 2286 -1995 2338
rect -1943 2286 -1923 2338
rect -1871 2286 -1851 2338
rect -1799 2286 -1779 2338
rect -1727 2286 -1707 2338
rect -1655 2286 -1635 2338
rect -1583 2286 -1563 2338
rect -1511 2286 -1491 2338
rect -1439 2286 -1419 2338
rect -1367 2286 -1347 2338
rect -1295 2286 -1275 2338
rect -1223 2286 -1203 2338
rect -1151 2286 -1131 2338
rect -1079 2286 -1059 2338
rect -1007 2286 -987 2338
rect -935 2286 -915 2338
rect -863 2286 -843 2338
rect -791 2286 -771 2338
rect -719 2286 -699 2338
rect -647 2286 -627 2338
rect -575 2286 -555 2338
rect -503 2286 -483 2338
rect -431 2286 -411 2338
rect -359 2286 -339 2338
rect -287 2286 -267 2338
rect -215 2286 -195 2338
rect -143 2286 -123 2338
rect -71 2286 -51 2338
rect 1 2286 21 2338
rect 73 2286 93 2338
rect 145 2286 165 2338
rect 217 2286 237 2338
rect 289 2286 309 2338
rect 361 2286 381 2338
rect 433 2286 453 2338
rect 505 2286 525 2338
rect 577 2286 597 2338
rect 649 2286 669 2338
rect 721 2286 741 2338
rect 793 2286 813 2338
rect 865 2286 885 2338
rect 937 2286 957 2338
rect 1009 2286 1029 2338
rect 1081 2286 1101 2338
rect 1153 2286 1173 2338
rect 1225 2286 1245 2338
rect 1297 2286 1317 2338
rect 1369 2286 1389 2338
rect 1441 2286 1461 2338
rect 1513 2286 1533 2338
rect 1585 2286 1605 2338
rect 1657 2286 1677 2338
rect 1729 2286 1749 2338
rect 1801 2286 1821 2338
rect 1873 2286 1893 2338
rect 1945 2286 1965 2338
rect 2017 2286 2037 2338
rect 2089 2286 2109 2338
rect 2161 2286 2181 2338
rect 2233 2286 2253 2338
rect 2305 2286 2325 2338
rect 2377 2286 2397 2338
rect 2449 2286 2469 2338
rect 2521 2286 2541 2338
rect 2593 2286 2613 2338
rect 2665 2286 2685 2338
rect 2737 2286 2757 2338
rect 2809 2286 2829 2338
rect 2881 2286 2901 2338
rect 2953 2286 2973 2338
rect 3025 2286 3045 2338
rect 3097 2286 3117 2338
rect 3169 2286 3189 2338
rect 3241 2286 3261 2338
rect 3313 2286 3333 2338
rect 3385 2286 3405 2338
rect 3457 2286 3477 2338
rect 3529 2286 3549 2338
rect 3601 2286 3621 2338
rect 3673 2286 3693 2338
rect 3745 2286 3765 2338
rect 3817 2286 3837 2338
rect 3889 2286 3909 2338
rect 3961 2286 3981 2338
rect 4033 2286 4039 2338
rect -3945 2266 4039 2286
rect -3945 2214 -3939 2266
rect -3887 2214 -3867 2266
rect -3815 2214 -3795 2266
rect -3743 2214 -3723 2266
rect -3671 2214 -3651 2266
rect -3599 2214 -3579 2266
rect -3527 2214 -3507 2266
rect -3455 2214 -3435 2266
rect -3383 2214 -3363 2266
rect -3311 2214 -3291 2266
rect -3239 2214 -3219 2266
rect -3167 2214 -3147 2266
rect -3095 2214 -3075 2266
rect -3023 2214 -3003 2266
rect -2951 2214 -2931 2266
rect -2879 2214 -2859 2266
rect -2807 2214 -2787 2266
rect -2735 2214 -2715 2266
rect -2663 2214 -2643 2266
rect -2591 2214 -2571 2266
rect -2519 2214 -2499 2266
rect -2447 2214 -2427 2266
rect -2375 2214 -2355 2266
rect -2303 2214 -2283 2266
rect -2231 2214 -2211 2266
rect -2159 2214 -2139 2266
rect -2087 2214 -2067 2266
rect -2015 2214 -1995 2266
rect -1943 2214 -1923 2266
rect -1871 2214 -1851 2266
rect -1799 2214 -1779 2266
rect -1727 2214 -1707 2266
rect -1655 2214 -1635 2266
rect -1583 2214 -1563 2266
rect -1511 2214 -1491 2266
rect -1439 2214 -1419 2266
rect -1367 2214 -1347 2266
rect -1295 2214 -1275 2266
rect -1223 2214 -1203 2266
rect -1151 2214 -1131 2266
rect -1079 2214 -1059 2266
rect -1007 2214 -987 2266
rect -935 2214 -915 2266
rect -863 2214 -843 2266
rect -791 2214 -771 2266
rect -719 2214 -699 2266
rect -647 2214 -627 2266
rect -575 2214 -555 2266
rect -503 2214 -483 2266
rect -431 2214 -411 2266
rect -359 2214 -339 2266
rect -287 2214 -267 2266
rect -215 2214 -195 2266
rect -143 2214 -123 2266
rect -71 2214 -51 2266
rect 1 2214 21 2266
rect 73 2214 93 2266
rect 145 2214 165 2266
rect 217 2214 237 2266
rect 289 2214 309 2266
rect 361 2214 381 2266
rect 433 2214 453 2266
rect 505 2214 525 2266
rect 577 2214 597 2266
rect 649 2214 669 2266
rect 721 2214 741 2266
rect 793 2214 813 2266
rect 865 2214 885 2266
rect 937 2214 957 2266
rect 1009 2214 1029 2266
rect 1081 2214 1101 2266
rect 1153 2214 1173 2266
rect 1225 2214 1245 2266
rect 1297 2214 1317 2266
rect 1369 2214 1389 2266
rect 1441 2214 1461 2266
rect 1513 2214 1533 2266
rect 1585 2214 1605 2266
rect 1657 2214 1677 2266
rect 1729 2214 1749 2266
rect 1801 2214 1821 2266
rect 1873 2214 1893 2266
rect 1945 2214 1965 2266
rect 2017 2214 2037 2266
rect 2089 2214 2109 2266
rect 2161 2214 2181 2266
rect 2233 2214 2253 2266
rect 2305 2214 2325 2266
rect 2377 2214 2397 2266
rect 2449 2214 2469 2266
rect 2521 2214 2541 2266
rect 2593 2214 2613 2266
rect 2665 2214 2685 2266
rect 2737 2214 2757 2266
rect 2809 2214 2829 2266
rect 2881 2214 2901 2266
rect 2953 2214 2973 2266
rect 3025 2214 3045 2266
rect 3097 2214 3117 2266
rect 3169 2214 3189 2266
rect 3241 2214 3261 2266
rect 3313 2214 3333 2266
rect 3385 2214 3405 2266
rect 3457 2214 3477 2266
rect 3529 2214 3549 2266
rect 3601 2214 3621 2266
rect 3673 2214 3693 2266
rect 3745 2214 3765 2266
rect 3817 2214 3837 2266
rect 3889 2214 3909 2266
rect 3961 2214 3981 2266
rect 4033 2214 4039 2266
rect -3945 2194 4039 2214
rect -3945 2142 -3939 2194
rect -3887 2142 -3867 2194
rect -3815 2142 -3795 2194
rect -3743 2142 -3723 2194
rect -3671 2142 -3651 2194
rect -3599 2142 -3579 2194
rect -3527 2142 -3507 2194
rect -3455 2142 -3435 2194
rect -3383 2142 -3363 2194
rect -3311 2142 -3291 2194
rect -3239 2142 -3219 2194
rect -3167 2142 -3147 2194
rect -3095 2142 -3075 2194
rect -3023 2142 -3003 2194
rect -2951 2142 -2931 2194
rect -2879 2142 -2859 2194
rect -2807 2142 -2787 2194
rect -2735 2142 -2715 2194
rect -2663 2142 -2643 2194
rect -2591 2142 -2571 2194
rect -2519 2142 -2499 2194
rect -2447 2142 -2427 2194
rect -2375 2142 -2355 2194
rect -2303 2142 -2283 2194
rect -2231 2142 -2211 2194
rect -2159 2142 -2139 2194
rect -2087 2142 -2067 2194
rect -2015 2142 -1995 2194
rect -1943 2142 -1923 2194
rect -1871 2142 -1851 2194
rect -1799 2142 -1779 2194
rect -1727 2142 -1707 2194
rect -1655 2142 -1635 2194
rect -1583 2142 -1563 2194
rect -1511 2142 -1491 2194
rect -1439 2142 -1419 2194
rect -1367 2142 -1347 2194
rect -1295 2142 -1275 2194
rect -1223 2142 -1203 2194
rect -1151 2142 -1131 2194
rect -1079 2142 -1059 2194
rect -1007 2142 -987 2194
rect -935 2142 -915 2194
rect -863 2142 -843 2194
rect -791 2142 -771 2194
rect -719 2142 -699 2194
rect -647 2142 -627 2194
rect -575 2142 -555 2194
rect -503 2142 -483 2194
rect -431 2142 -411 2194
rect -359 2142 -339 2194
rect -287 2142 -267 2194
rect -215 2142 -195 2194
rect -143 2142 -123 2194
rect -71 2142 -51 2194
rect 1 2142 21 2194
rect 73 2142 93 2194
rect 145 2142 165 2194
rect 217 2142 237 2194
rect 289 2142 309 2194
rect 361 2142 381 2194
rect 433 2142 453 2194
rect 505 2142 525 2194
rect 577 2142 597 2194
rect 649 2142 669 2194
rect 721 2142 741 2194
rect 793 2142 813 2194
rect 865 2142 885 2194
rect 937 2142 957 2194
rect 1009 2142 1029 2194
rect 1081 2142 1101 2194
rect 1153 2142 1173 2194
rect 1225 2142 1245 2194
rect 1297 2142 1317 2194
rect 1369 2142 1389 2194
rect 1441 2142 1461 2194
rect 1513 2142 1533 2194
rect 1585 2142 1605 2194
rect 1657 2142 1677 2194
rect 1729 2142 1749 2194
rect 1801 2142 1821 2194
rect 1873 2142 1893 2194
rect 1945 2142 1965 2194
rect 2017 2142 2037 2194
rect 2089 2142 2109 2194
rect 2161 2142 2181 2194
rect 2233 2142 2253 2194
rect 2305 2142 2325 2194
rect 2377 2142 2397 2194
rect 2449 2142 2469 2194
rect 2521 2142 2541 2194
rect 2593 2142 2613 2194
rect 2665 2142 2685 2194
rect 2737 2142 2757 2194
rect 2809 2142 2829 2194
rect 2881 2142 2901 2194
rect 2953 2142 2973 2194
rect 3025 2142 3045 2194
rect 3097 2142 3117 2194
rect 3169 2142 3189 2194
rect 3241 2142 3261 2194
rect 3313 2142 3333 2194
rect 3385 2142 3405 2194
rect 3457 2142 3477 2194
rect 3529 2142 3549 2194
rect 3601 2142 3621 2194
rect 3673 2142 3693 2194
rect 3745 2142 3765 2194
rect 3817 2142 3837 2194
rect 3889 2142 3909 2194
rect 3961 2142 3981 2194
rect 4033 2142 4039 2194
rect -3945 2136 4039 2142
rect -3938 4 -3800 10
rect -3938 -48 -3932 4
rect -3880 -48 -3858 4
rect -3806 -48 -3800 4
rect -3938 -70 -3800 -48
rect -3938 -122 -3932 -70
rect -3880 -122 -3858 -70
rect -3806 -122 -3800 -70
rect -3938 -128 -3800 -122
use nfet$10  nfet$10_0
timestamp 1698900908
transform 0 -1 2047 1 0 149
box -26 -40 690 6106
use nfet  nfet_0
timestamp 1698900908
transform 0 -1 -3769 -1 0 117
box -26 -40 276 306
use pfet$6  pfet$6_0
timestamp 1698900908
transform 0 -1 4047 1 0 899
box -61 -76 1534 8144
<< labels >>
flabel metal1 s -4099 -20 -3983 92 0 FreeSans 44 0 0 0 CTRL
port 2 nsew
flabel metal1 s -3942 688 4036 1096 0 FreeSans 44 0 0 0 OUT
port 3 nsew
flabel metal1 s -3852 909 -3852 909 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 178 907 178 907 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 2245 914 2245 914 0 FreeSans 44 0 0 0 OUT
flabel metal1 s -2064 943 -2064 943 0 FreeSans 44 0 0 0 OUT
flabel metal1 s -4118 308 -4003 1892 0 FreeSans 44 0 0 0 IN
port 4 nsew
flabel metal1 s -4063 333 -4063 333 0 FreeSans 44 0 0 0 IN
flabel metal1 s -4062 1220 -4062 1220 0 FreeSans 44 0 0 0 IN
flabel metal1 s -4062 1587 -4062 1587 0 FreeSans 44 0 0 0 IN
flabel metal1 s -4060 834 -4060 834 0 FreeSans 44 0 0 0 IN
flabel metal2 s -3938 -128 -3800 10 0 FreeSans 44 0 0 0 VSS
port 6 nsew
flabel metal2 s -3945 2135 4039 2343 0 FreeSans 44 0 0 0 VDD
port 7 nsew
flabel metal2 s 3994 2243 3994 2243 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 9 2237 9 2237 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 2352 2229 2352 2229 0 FreeSans 44 0 0 0 VDD
flabel metal2 s -2016 2250 -2016 2250 0 FreeSans 44 0 0 0 VDD
<< end >>
