magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< xpolycontact >>
rect -35 46 35 482
rect -35 -482 35 -46
<< ppolyres >>
rect -35 -46 35 46
<< viali >>
rect -17 429 17 463
rect -17 357 17 391
rect -17 285 17 319
rect -17 213 17 247
rect -17 141 17 175
rect -17 69 17 103
rect -17 -102 17 -68
rect -17 -174 17 -140
rect -17 -246 17 -212
rect -17 -318 17 -284
rect -17 -390 17 -356
rect -17 -462 17 -428
<< metal1 >>
rect -25 463 25 476
rect -25 429 -17 463
rect 17 429 25 463
rect -25 391 25 429
rect -25 357 -17 391
rect 17 357 25 391
rect -25 319 25 357
rect -25 285 -17 319
rect 17 285 25 319
rect -25 247 25 285
rect -25 213 -17 247
rect 17 213 25 247
rect -25 175 25 213
rect -25 141 -17 175
rect 17 141 25 175
rect -25 103 25 141
rect -25 69 -17 103
rect 17 69 25 103
rect -25 55 25 69
rect -25 -68 25 -55
rect -25 -102 -17 -68
rect 17 -102 25 -68
rect -25 -140 25 -102
rect -25 -174 -17 -140
rect 17 -174 25 -140
rect -25 -212 25 -174
rect -25 -246 -17 -212
rect 17 -246 25 -212
rect -25 -284 25 -246
rect -25 -318 -17 -284
rect 17 -318 25 -284
rect -25 -356 25 -318
rect -25 -390 -17 -356
rect 17 -390 25 -356
rect -25 -428 25 -390
rect -25 -462 -17 -428
rect 17 -462 25 -428
rect -25 -476 25 -462
<< end >>
