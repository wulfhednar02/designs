magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -635 -2610 635 2610
<< l66d20 >>
rect -175 -2410 175 2410
<< l94d20 >>
rect -285 -2520 285 2520
<< l86d20 >>
rect -635 -2610 635 2610
<< l66d44 >>
rect -95 330 95 2330
rect -95 -2330 95 -330
<< l67d44 >>
rect -85 345 85 515
rect -85 705 85 875
rect -85 1065 85 1235
rect -85 1425 85 1595
rect -85 1785 85 1955
rect -85 2145 85 2315
rect -85 -2310 85 -2140
rect -85 -1950 85 -1780
rect -85 -1590 85 -1420
rect -85 -1230 85 -1060
rect -85 -870 85 -700
rect -85 -510 85 -340
<< l95d20 >>
rect -270 -2505 270 2505
<< l67d20 >>
rect -175 250 175 2410
rect -175 -2410 175 -250
<< l66d13 >>
rect -175 -310 175 310
<< l68d20 >>
rect -125 276 125 2380
rect -125 -2380 125 -276
<< end >>
