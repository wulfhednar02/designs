magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< error_s >>
rect 44541 40557 44553 40563
rect 44563 40557 44575 40563
rect 44529 40539 44530 40551
rect 44585 40539 44587 40551
rect 41271 40413 41277 40419
rect 41301 40389 41307 40409
rect 41343 40301 41349 40321
rect 41301 40279 41307 40285
rect 44529 40171 44530 40183
rect 44585 40171 44587 40183
rect 44541 40159 44553 40165
rect 44563 40159 44575 40165
<< locali >>
rect 41155 40341 41219 40360
rect 41155 40307 41163 40341
rect 41197 40307 41219 40341
rect 41155 40286 41219 40307
rect 41457 40304 41502 40344
rect 42383 40304 42595 40344
<< viali >>
rect 44447 40616 44481 40650
rect 44539 40616 44573 40650
rect 44541 40517 44575 40551
rect 44541 40431 44575 40465
rect 44541 40344 44575 40378
rect 41163 40307 41197 40341
rect 41242 40307 41276 40341
rect 44541 40257 44575 40291
rect 44541 40171 44575 40205
rect 44447 40072 44481 40106
rect 44539 40072 44573 40106
<< metal1 >>
rect 44530 40551 44585 40557
rect 44530 40517 44541 40551
rect 44575 40517 44585 40551
rect 44530 40465 44585 40517
rect 44530 40431 44541 40465
rect 44575 40431 44585 40465
rect 44530 40378 44585 40431
rect 41155 40341 41287 40360
rect 41155 40307 41163 40341
rect 41197 40307 41242 40341
rect 41276 40307 41287 40341
rect 41155 40286 41287 40307
rect 44530 40344 44541 40378
rect 44575 40344 44585 40378
rect 44530 40291 44585 40344
rect 44530 40257 44541 40291
rect 44575 40257 44585 40291
rect 44530 40205 44585 40257
rect 44530 40171 44541 40205
rect 44575 40171 44585 40205
rect 44530 40165 44585 40171
<< via1 >>
rect 41218 40607 41270 40659
rect 41310 40607 41362 40659
rect 41402 40607 41454 40659
rect 41494 40607 41546 40659
rect 41586 40607 41638 40659
rect 41678 40607 41730 40659
rect 41770 40607 41822 40659
rect 41862 40607 41914 40659
rect 41954 40607 42006 40659
rect 42046 40607 42098 40659
rect 42138 40607 42190 40659
rect 42230 40607 42282 40659
rect 42322 40607 42374 40659
rect 42414 40607 42466 40659
rect 42506 40607 42558 40659
rect 42598 40607 42650 40659
rect 42690 40607 42742 40659
rect 42782 40607 42834 40659
rect 42874 40607 42926 40659
rect 42966 40607 43018 40659
rect 43058 40607 43110 40659
rect 43150 40607 43202 40659
rect 43242 40607 43294 40659
rect 43334 40607 43386 40659
rect 43426 40607 43478 40659
rect 43518 40607 43570 40659
rect 43610 40607 43662 40659
rect 43702 40607 43754 40659
rect 43794 40607 43846 40659
rect 43886 40607 43938 40659
rect 43978 40607 44030 40659
rect 44070 40607 44122 40659
rect 44162 40607 44214 40659
rect 44254 40607 44306 40659
rect 44346 40607 44398 40659
rect 44438 40650 44490 40659
rect 44438 40616 44447 40650
rect 44447 40616 44481 40650
rect 44481 40616 44490 40650
rect 44438 40607 44490 40616
rect 44530 40650 44582 40659
rect 44530 40616 44539 40650
rect 44539 40616 44573 40650
rect 44573 40616 44582 40650
rect 44530 40607 44582 40616
rect 41218 40063 41270 40115
rect 41310 40063 41362 40115
rect 41402 40063 41454 40115
rect 41494 40063 41546 40115
rect 41586 40063 41638 40115
rect 41678 40063 41730 40115
rect 41770 40063 41822 40115
rect 41862 40063 41914 40115
rect 41954 40063 42006 40115
rect 42046 40063 42098 40115
rect 42138 40063 42190 40115
rect 42230 40063 42282 40115
rect 42322 40063 42374 40115
rect 42414 40063 42466 40115
rect 42506 40063 42558 40115
rect 42598 40063 42650 40115
rect 42690 40063 42742 40115
rect 42782 40063 42834 40115
rect 42874 40063 42926 40115
rect 42966 40063 43018 40115
rect 43058 40063 43110 40115
rect 43150 40063 43202 40115
rect 43242 40063 43294 40115
rect 43334 40063 43386 40115
rect 43426 40063 43478 40115
rect 43518 40063 43570 40115
rect 43610 40063 43662 40115
rect 43702 40063 43754 40115
rect 43794 40063 43846 40115
rect 43886 40063 43938 40115
rect 43978 40063 44030 40115
rect 44070 40063 44122 40115
rect 44162 40063 44214 40115
rect 44254 40063 44306 40115
rect 44346 40063 44398 40115
rect 44438 40106 44490 40115
rect 44438 40072 44447 40106
rect 44447 40072 44481 40106
rect 44481 40072 44490 40106
rect 44438 40063 44490 40072
rect 44530 40106 44582 40115
rect 44530 40072 44539 40106
rect 44539 40072 44573 40106
rect 44573 40072 44582 40106
rect 44530 40063 44582 40072
<< metal2 >>
rect 41198 40659 44602 40681
rect 41198 40607 41218 40659
rect 41270 40607 41310 40659
rect 41362 40607 41402 40659
rect 41454 40607 41494 40659
rect 41546 40607 41586 40659
rect 41638 40607 41678 40659
rect 41730 40607 41770 40659
rect 41822 40607 41862 40659
rect 41914 40607 41954 40659
rect 42006 40607 42046 40659
rect 42098 40607 42138 40659
rect 42190 40607 42230 40659
rect 42282 40607 42322 40659
rect 42374 40607 42414 40659
rect 42466 40607 42506 40659
rect 42558 40607 42598 40659
rect 42650 40607 42690 40659
rect 42742 40607 42782 40659
rect 42834 40607 42874 40659
rect 42926 40607 42966 40659
rect 43018 40607 43058 40659
rect 43110 40607 43150 40659
rect 43202 40607 43242 40659
rect 43294 40607 43334 40659
rect 43386 40607 43426 40659
rect 43478 40607 43518 40659
rect 43570 40607 43610 40659
rect 43662 40607 43702 40659
rect 43754 40607 43794 40659
rect 43846 40607 43886 40659
rect 43938 40607 43978 40659
rect 44030 40607 44070 40659
rect 44122 40607 44162 40659
rect 44214 40607 44254 40659
rect 44306 40607 44346 40659
rect 44398 40607 44438 40659
rect 44490 40607 44530 40659
rect 44582 40607 44602 40659
rect 41198 40585 44602 40607
rect 41198 40115 44602 40137
rect 41198 40063 41218 40115
rect 41270 40063 41310 40115
rect 41362 40063 41402 40115
rect 41454 40063 41494 40115
rect 41546 40063 41586 40115
rect 41638 40063 41678 40115
rect 41730 40063 41770 40115
rect 41822 40063 41862 40115
rect 41914 40063 41954 40115
rect 42006 40063 42046 40115
rect 42098 40063 42138 40115
rect 42190 40063 42230 40115
rect 42282 40063 42322 40115
rect 42374 40063 42414 40115
rect 42466 40063 42506 40115
rect 42558 40063 42598 40115
rect 42650 40063 42690 40115
rect 42742 40063 42782 40115
rect 42834 40063 42874 40115
rect 42926 40063 42966 40115
rect 43018 40063 43058 40115
rect 43110 40063 43150 40115
rect 43202 40063 43242 40115
rect 43294 40063 43334 40115
rect 43386 40063 43426 40115
rect 43478 40063 43518 40115
rect 43570 40063 43610 40115
rect 43662 40063 43702 40115
rect 43754 40063 43794 40115
rect 43846 40063 43886 40115
rect 43938 40063 43978 40115
rect 44030 40063 44070 40115
rect 44122 40063 44162 40115
rect 44214 40063 44254 40115
rect 44306 40063 44346 40115
rect 44398 40063 44438 40115
rect 44490 40063 44530 40115
rect 44582 40063 44602 40115
rect 41198 40041 44602 40063
use sky130_fd_sc_hd__buf_1  sky130_fd_sc_hd__buf_1_0
timestamp 1698900908
transform 1 0 41198 0 1 40089
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  sky130_fd_sc_hd__buf_8_0
timestamp 1698900908
transform 1 0 41474 0 1 40089
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_16  sky130_fd_sc_hd__buf_16_0
timestamp 1698900908
transform 1 0 42578 0 1 40089
box -38 -48 2062 592
<< labels >>
flabel metal1 s 41155 40286 41287 40360 0 FreeSans 44 0 0 0 IN
port 2 nsew
flabel metal1 s 44530 40167 44585 40556 0 FreeSans 44 0 0 0 OUT
port 3 nsew
flabel metal1 s 44557 40183 44557 40183 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 44558 40361 44558 40361 0 FreeSans 44 0 0 0 OUT
flabel metal2 s 41198 40041 44602 40137 0 FreeSans 44 0 0 0 VSS
port 5 nsew
flabel metal2 s 44564 40091 44564 40091 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 42890 40094 42890 40094 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 41942 40091 41942 40091 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 43811 40098 43811 40098 0 FreeSans 44 0 0 0 VSS
flabel metal2 s 41198 40585 44602 40681 0 FreeSans 44 0 0 0 VDD
port 6 nsew
flabel metal2 s 44551 40639 44551 40639 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 42887 40637 42887 40637 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 41951 40635 41951 40635 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 43830 40637 43830 40637 0 FreeSans 44 0 0 0 VDD
<< end >>
