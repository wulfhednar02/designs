magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -20590 -789 20615 12166
<< l67d44 >>
rect 150 10753 320 10923
rect 150 11113 320 11283
rect 150 11473 320 11643
rect 10230 10753 10400 10923
rect 10590 10753 10760 10923
rect 10950 10753 11120 10923
rect 11310 10753 11480 10923
rect 11670 10753 11840 10923
rect 12030 10753 12200 10923
rect 12390 10753 12560 10923
rect 12750 10753 12920 10923
rect 13110 10753 13280 10923
rect 13470 10753 13640 10923
rect 13830 10753 14000 10923
rect 14190 10753 14360 10923
rect 14550 10753 14720 10923
rect 14910 10753 15080 10923
rect 15270 10753 15440 10923
rect 15630 10753 15800 10923
rect 15990 10753 16160 10923
rect 16350 10753 16520 10923
rect 16710 10753 16880 10923
rect 17070 10753 17240 10923
rect 17430 10753 17600 10923
rect 17790 10753 17960 10923
rect 18150 10753 18320 10923
rect 18510 10753 18680 10923
rect 18870 10753 19040 10923
rect 19230 10753 19400 10923
rect 19590 10753 19760 10923
rect 19950 10753 20120 10923
rect 10230 11113 10400 11283
rect 10590 11113 10760 11283
rect 10950 11113 11120 11283
rect 11310 11113 11480 11283
rect 11670 11113 11840 11283
rect 12030 11113 12200 11283
rect 12390 11113 12560 11283
rect 12750 11113 12920 11283
rect 13110 11113 13280 11283
rect 13470 11113 13640 11283
rect 13830 11113 14000 11283
rect 14190 11113 14360 11283
rect 14550 11113 14720 11283
rect 14910 11113 15080 11283
rect 15270 11113 15440 11283
rect 15630 11113 15800 11283
rect 15990 11113 16160 11283
rect 16350 11113 16520 11283
rect 16710 11113 16880 11283
rect 17070 11113 17240 11283
rect 17430 11113 17600 11283
rect 17790 11113 17960 11283
rect 18150 11113 18320 11283
rect 18510 11113 18680 11283
rect 18870 11113 19040 11283
rect 19230 11113 19400 11283
rect 19590 11113 19760 11283
rect 19950 11113 20120 11283
rect 10230 11473 10400 11643
rect 10590 11473 10760 11643
rect 10950 11473 11120 11643
rect 11310 11473 11480 11643
rect 11670 11473 11840 11643
rect 12030 11473 12200 11643
rect 12390 11473 12560 11643
rect 12750 11473 12920 11643
rect 13110 11473 13280 11643
rect 13470 11473 13640 11643
rect 13830 11473 14000 11643
rect 14190 11473 14360 11643
rect 14550 11473 14720 11643
rect 14910 11473 15080 11643
rect 15270 11473 15440 11643
rect 15630 11473 15800 11643
rect 15990 11473 16160 11643
rect 16350 11473 16520 11643
rect 16710 11473 16880 11643
rect 17070 11473 17240 11643
rect 17430 11473 17600 11643
rect 17790 11473 17960 11643
rect 18150 11473 18320 11643
rect 18510 11473 18680 11643
rect 18870 11473 19040 11643
rect 19230 11473 19400 11643
rect 19590 11473 19760 11643
rect 19950 11473 20120 11643
rect 3390 10753 3560 10923
rect 3750 10753 3920 10923
rect 4110 10753 4280 10923
rect 4470 10753 4640 10923
rect 4830 10753 5000 10923
rect 5190 10753 5360 10923
rect 5550 10753 5720 10923
rect 5910 10753 6080 10923
rect 6270 10753 6440 10923
rect 6630 10753 6800 10923
rect 6990 10753 7160 10923
rect 7350 10753 7520 10923
rect 7710 10753 7880 10923
rect 8070 10753 8240 10923
rect 8430 10753 8600 10923
rect 8790 10753 8960 10923
rect 9150 10753 9320 10923
rect 9510 10753 9680 10923
rect 9870 10753 10040 10923
rect 1230 10753 1400 10923
rect 1590 10753 1760 10923
rect 1950 10753 2120 10923
rect 510 10753 680 10923
rect 510 11113 680 11283
rect 870 11113 1040 11283
rect 870 10753 1040 10923
rect 510 11473 680 11643
rect 870 11473 1040 11643
rect 1230 11473 1400 11643
rect 1590 11473 1760 11643
rect 1950 11473 2120 11643
rect 2310 11473 2480 11643
rect 2670 11473 2840 11643
rect 3030 11473 3200 11643
rect 3390 11473 3560 11643
rect 3750 11473 3920 11643
rect 4110 11473 4280 11643
rect 4470 11473 4640 11643
rect 4830 11473 5000 11643
rect 5190 11473 5360 11643
rect 5550 11473 5720 11643
rect 5910 11473 6080 11643
rect 6270 11473 6440 11643
rect 6630 11473 6800 11643
rect 6990 11473 7160 11643
rect 7350 11473 7520 11643
rect 7710 11473 7880 11643
rect 8070 11473 8240 11643
rect 8430 11473 8600 11643
rect 8790 11473 8960 11643
rect 9150 11473 9320 11643
rect 9510 11473 9680 11643
rect 9870 11473 10040 11643
rect 1230 11113 1400 11283
rect 1590 11113 1760 11283
rect 1950 11113 2120 11283
rect 2310 11113 2480 11283
rect 2670 11113 2840 11283
rect 3030 11113 3200 11283
rect 3390 11113 3560 11283
rect 3750 11113 3920 11283
rect 4110 11113 4280 11283
rect 4470 11113 4640 11283
rect 4830 11113 5000 11283
rect 5190 11113 5360 11283
rect 5550 11113 5720 11283
rect 5910 11113 6080 11283
rect 6270 11113 6440 11283
rect 6630 11113 6800 11283
rect 6990 11113 7160 11283
rect 7350 11113 7520 11283
rect 7710 11113 7880 11283
rect 8070 11113 8240 11283
rect 8430 11113 8600 11283
rect 8790 11113 8960 11283
rect 9150 11113 9320 11283
rect 9510 11113 9680 11283
rect 9870 11113 10040 11283
rect 2310 10753 2480 10923
rect 2670 10753 2840 10923
rect 3030 10753 3200 10923
rect -9570 11113 -9400 11283
rect -9210 11113 -9040 11283
rect -8850 11113 -8680 11283
rect -8490 11113 -8320 11283
rect -8130 11113 -7960 11283
rect -7770 11113 -7600 11283
rect -7410 11113 -7240 11283
rect -7050 11113 -6880 11283
rect -6690 11113 -6520 11283
rect -6330 11113 -6160 11283
rect -5970 11113 -5800 11283
rect -5610 11113 -5440 11283
rect -5250 11113 -5080 11283
rect -4890 11113 -4720 11283
rect -4530 11113 -4360 11283
rect -4170 11113 -4000 11283
rect -3810 11113 -3640 11283
rect -3450 11113 -3280 11283
rect -3090 11113 -2920 11283
rect -2730 11113 -2560 11283
rect -2370 11113 -2200 11283
rect -2010 11113 -1840 11283
rect -1650 11113 -1480 11283
rect -1290 11113 -1120 11283
rect -930 11113 -760 11283
rect -570 11113 -400 11283
rect -210 11113 -40 11283
rect -9570 10753 -9400 10923
rect -9210 10753 -9040 10923
rect -8850 10753 -8680 10923
rect -8490 10753 -8320 10923
rect -8130 10753 -7960 10923
rect -7770 10753 -7600 10923
rect -7410 10753 -7240 10923
rect -7050 10753 -6880 10923
rect -6690 10753 -6520 10923
rect -6330 10753 -6160 10923
rect -5970 10753 -5800 10923
rect -5610 10753 -5440 10923
rect -5250 10753 -5080 10923
rect -4890 10753 -4720 10923
rect -4530 10753 -4360 10923
rect -4170 10753 -4000 10923
rect -3810 10753 -3640 10923
rect -3450 10753 -3280 10923
rect -3090 10753 -2920 10923
rect -2730 10753 -2560 10923
rect -2370 10753 -2200 10923
rect -2010 10753 -1840 10923
rect -1650 10753 -1480 10923
rect -1290 10753 -1120 10923
rect -930 10753 -760 10923
rect -570 10753 -400 10923
rect -210 10753 -40 10923
rect -9570 11473 -9400 11643
rect -9210 11473 -9040 11643
rect -8850 11473 -8680 11643
rect -8490 11473 -8320 11643
rect -8130 11473 -7960 11643
rect -7770 11473 -7600 11643
rect -7410 11473 -7240 11643
rect -7050 11473 -6880 11643
rect -6690 11473 -6520 11643
rect -6330 11473 -6160 11643
rect -5970 11473 -5800 11643
rect -5610 11473 -5440 11643
rect -5250 11473 -5080 11643
rect -4890 11473 -4720 11643
rect -4530 11473 -4360 11643
rect -4170 11473 -4000 11643
rect -3810 11473 -3640 11643
rect -3450 11473 -3280 11643
rect -3090 11473 -2920 11643
rect -2730 11473 -2560 11643
rect -2370 11473 -2200 11643
rect -2010 11473 -1840 11643
rect -1650 11473 -1480 11643
rect -1290 11473 -1120 11643
rect -930 11473 -760 11643
rect -570 11473 -400 11643
rect -210 11473 -40 11643
rect -17850 11113 -17680 11283
rect -17490 11113 -17320 11283
rect -17130 11113 -16960 11283
rect -16770 11113 -16600 11283
rect -16410 11113 -16240 11283
rect -16050 11113 -15880 11283
rect -15690 11113 -15520 11283
rect -15330 11113 -15160 11283
rect -14970 11113 -14800 11283
rect -14610 11113 -14440 11283
rect -14250 11113 -14080 11283
rect -13890 11113 -13720 11283
rect -13530 11113 -13360 11283
rect -13170 11113 -13000 11283
rect -12810 11113 -12640 11283
rect -12450 11113 -12280 11283
rect -12090 11113 -11920 11283
rect -11730 11113 -11560 11283
rect -11370 11113 -11200 11283
rect -11010 11113 -10840 11283
rect -10650 11113 -10480 11283
rect -10290 11113 -10120 11283
rect -9930 11113 -9760 11283
rect -18930 11113 -18760 11283
rect -18930 10753 -18760 10923
rect -19650 10753 -19480 10923
rect -19290 10753 -19120 10923
rect -19290 11113 -19120 11283
rect -19290 11473 -19120 11643
rect -18930 11473 -18760 11643
rect -18570 11473 -18400 11643
rect -18210 11473 -18040 11643
rect -17850 11473 -17680 11643
rect -17490 11473 -17320 11643
rect -17130 11473 -16960 11643
rect -16770 11473 -16600 11643
rect -16410 11473 -16240 11643
rect -16050 11473 -15880 11643
rect -15690 11473 -15520 11643
rect -15330 11473 -15160 11643
rect -14970 11473 -14800 11643
rect -14610 11473 -14440 11643
rect -14250 11473 -14080 11643
rect -13890 11473 -13720 11643
rect -13530 11473 -13360 11643
rect -13170 11473 -13000 11643
rect -12810 11473 -12640 11643
rect -12450 11473 -12280 11643
rect -12090 11473 -11920 11643
rect -11730 11473 -11560 11643
rect -11370 11473 -11200 11643
rect -11010 11473 -10840 11643
rect -10650 11473 -10480 11643
rect -10290 11473 -10120 11643
rect -9930 11473 -9760 11643
rect -18570 10753 -18400 10923
rect -18210 10753 -18040 10923
rect -17850 10753 -17680 10923
rect -17490 10753 -17320 10923
rect -17130 10753 -16960 10923
rect -16770 10753 -16600 10923
rect -16410 10753 -16240 10923
rect -16050 10753 -15880 10923
rect -15690 10753 -15520 10923
rect -15330 10753 -15160 10923
rect -14970 10753 -14800 10923
rect -14610 10753 -14440 10923
rect -14250 10753 -14080 10923
rect -13890 10753 -13720 10923
rect -13530 10753 -13360 10923
rect -13170 10753 -13000 10923
rect -12810 10753 -12640 10923
rect -12450 10753 -12280 10923
rect -12090 10753 -11920 10923
rect -11730 10753 -11560 10923
rect -11370 10753 -11200 10923
rect -11010 10753 -10840 10923
rect -10650 10753 -10480 10923
rect -10290 10753 -10120 10923
rect -9930 10753 -9760 10923
rect -18570 11113 -18400 11283
rect -18210 11113 -18040 11283
rect -19650 11113 -19480 11283
rect -19650 11473 -19480 11643
rect -19250 -525 -19080 -355
rect -19610 -525 -19440 -355
<< l68d20 >>
rect -20245 3270 -20015 5570
rect -19690 -640 -19000 50
rect -19710 3440 20180 5480
rect -20551 -157 -19871 523
rect -20590 1540 -20015 9460
rect -19710 3440 20180 5480
rect -20590 1540 -20015 9460
rect -19690 320 -19000 1370
rect -19710 10500 20180 11688
rect 20180 10753 20200 11688
rect -19730 10753 -19710 11688
<< l68d16 >>
rect -19710 3440 20180 5480
rect -20590 1540 -20015 9460
rect -20496 -102 -19916 463
<< l68d44 >>
rect 160 10763 310 10913
rect 160 11123 310 11273
rect 160 11483 310 11633
rect 12400 11123 12550 11273
rect 12760 11123 12910 11273
rect 13120 11123 13270 11273
rect 17080 11483 17230 11633
rect 13480 11123 13630 11273
rect 17440 11483 17590 11633
rect 13840 11123 13990 11273
rect 17800 11483 17950 11633
rect 14200 11123 14350 11273
rect 18160 11483 18310 11633
rect 14560 11123 14710 11273
rect 18520 11483 18670 11633
rect 14920 11123 15070 11273
rect 18880 11483 19030 11633
rect 15280 11123 15430 11273
rect 19240 11483 19390 11633
rect 15640 11123 15790 11273
rect 19600 11483 19750 11633
rect 16000 11123 16150 11273
rect 19960 11483 20110 11633
rect 16360 11123 16510 11273
rect 10240 10763 10390 10913
rect 16720 11123 16870 11273
rect 10600 10763 10750 10913
rect 17080 11123 17230 11273
rect 10960 10763 11110 10913
rect 17440 11123 17590 11273
rect 11320 10763 11470 10913
rect 17800 11123 17950 11273
rect 11680 10763 11830 10913
rect 18160 11123 18310 11273
rect 12040 10763 12190 10913
rect 18520 11123 18670 11273
rect 12400 10763 12550 10913
rect 18880 11123 19030 11273
rect 12760 10763 12910 10913
rect 19240 11123 19390 11273
rect 13120 10763 13270 10913
rect 19600 11123 19750 11273
rect 13480 10763 13630 10913
rect 19960 11123 20110 11273
rect 13840 10763 13990 10913
rect 10240 11483 10390 11633
rect 14200 10763 14350 10913
rect 10600 11483 10750 11633
rect 14560 10763 14710 10913
rect 10960 11483 11110 11633
rect 14920 10763 15070 10913
rect 11320 11483 11470 11633
rect 15280 10763 15430 10913
rect 11680 11483 11830 11633
rect 15640 10763 15790 10913
rect 12040 11483 12190 11633
rect 16000 10763 16150 10913
rect 12400 11483 12550 11633
rect 12760 11483 12910 11633
rect 16360 10763 16510 10913
rect 13120 11483 13270 11633
rect 16720 10763 16870 10913
rect 17080 10763 17230 10913
rect 13480 11483 13630 11633
rect 17440 10763 17590 10913
rect 17800 10763 17950 10913
rect 13840 11483 13990 11633
rect 18160 10763 18310 10913
rect 18520 10763 18670 10913
rect 14200 11483 14350 11633
rect 18880 10763 19030 10913
rect 19240 10763 19390 10913
rect 14560 11483 14710 11633
rect 19600 10763 19750 10913
rect 19960 10763 20110 10913
rect 14920 11483 15070 11633
rect 15280 11483 15430 11633
rect 15640 11483 15790 11633
rect 16000 11483 16150 11633
rect 16360 11483 16510 11633
rect 16720 11483 16870 11633
rect 10240 11123 10390 11273
rect 10600 11123 10750 11273
rect 10960 11123 11110 11273
rect 11320 11123 11470 11273
rect 11680 11123 11830 11273
rect 12040 11123 12190 11273
rect 2320 11123 2470 11273
rect 2680 11123 2830 11273
rect 3040 11123 3190 11273
rect 3400 11123 3550 11273
rect 3760 11123 3910 11273
rect 4120 11123 4270 11273
rect 4480 11123 4630 11273
rect 4840 11123 4990 11273
rect 5200 11123 5350 11273
rect 1240 11123 1390 11273
rect 1600 11123 1750 11273
rect 1960 11123 2110 11273
rect 9880 10763 10030 10913
rect 9880 11483 10030 11633
rect 880 11483 1030 11633
rect 3040 11483 3190 11633
rect 3400 11483 3550 11633
rect 1240 11483 1390 11633
rect 3760 11483 3910 11633
rect 4120 11483 4270 11633
rect 1600 11483 1750 11633
rect 4480 11483 4630 11633
rect 4840 11483 4990 11633
rect 1960 11483 2110 11633
rect 5200 11483 5350 11633
rect 5560 11483 5710 11633
rect 2320 11483 2470 11633
rect 5920 11483 6070 11633
rect 6280 11483 6430 11633
rect 2680 11483 2830 11633
rect 5920 11123 6070 11273
rect 520 10763 670 10913
rect 880 10763 1030 10913
rect 1240 10763 1390 10913
rect 1600 10763 1750 10913
rect 1960 10763 2110 10913
rect 2320 10763 2470 10913
rect 2680 10763 2830 10913
rect 3040 10763 3190 10913
rect 3400 10763 3550 10913
rect 3760 10763 3910 10913
rect 4120 10763 4270 10913
rect 4480 10763 4630 10913
rect 4840 10763 4990 10913
rect 5200 10763 5350 10913
rect 5560 10763 5710 10913
rect 5920 10763 6070 10913
rect 6280 10763 6430 10913
rect 6640 10763 6790 10913
rect 7000 10763 7150 10913
rect 7360 10763 7510 10913
rect 7720 10763 7870 10913
rect 8080 10763 8230 10913
rect 8440 10763 8590 10913
rect 8800 10763 8950 10913
rect 9160 10763 9310 10913
rect 9520 10763 9670 10913
rect 6280 11123 6430 11273
rect 6640 11483 6790 11633
rect 7000 11483 7150 11633
rect 7360 11483 7510 11633
rect 7720 11483 7870 11633
rect 8080 11483 8230 11633
rect 8440 11483 8590 11633
rect 8800 11483 8950 11633
rect 9160 11483 9310 11633
rect 9520 11483 9670 11633
rect 520 11123 670 11273
rect 9520 11123 9670 11273
rect 880 11123 1030 11273
rect 6640 11123 6790 11273
rect 7000 11123 7150 11273
rect 7360 11123 7510 11273
rect 7720 11123 7870 11273
rect 8080 11123 8230 11273
rect 8440 11123 8590 11273
rect 8800 11123 8950 11273
rect 9160 11123 9310 11273
rect 5560 11123 5710 11273
rect 520 11483 670 11633
rect 9880 11123 10030 11273
rect -200 11123 -50 11273
rect -200 10763 -50 10913
rect -200 11483 -50 11633
rect -7400 11483 -7250 11633
rect -7040 11483 -6890 11633
rect -6680 11483 -6530 11633
rect -6320 11483 -6170 11633
rect -5960 11483 -5810 11633
rect -5600 11483 -5450 11633
rect -5240 11483 -5090 11633
rect -4880 11483 -4730 11633
rect -4520 11483 -4370 11633
rect -4160 11483 -4010 11633
rect -3800 11483 -3650 11633
rect -3440 11483 -3290 11633
rect -3080 11483 -2930 11633
rect -2720 11483 -2570 11633
rect -2360 11483 -2210 11633
rect -2000 11483 -1850 11633
rect -1640 11483 -1490 11633
rect -1280 11483 -1130 11633
rect -920 11483 -770 11633
rect -560 11483 -410 11633
rect -9200 10763 -9050 10913
rect -9560 11123 -9410 11273
rect -9200 11123 -9050 11273
rect -8840 11123 -8690 11273
rect -8480 11123 -8330 11273
rect -8120 11123 -7970 11273
rect -7760 11123 -7610 11273
rect -7400 11123 -7250 11273
rect -7040 11123 -6890 11273
rect -6680 11123 -6530 11273
rect -6320 11123 -6170 11273
rect -5960 11123 -5810 11273
rect -5600 11123 -5450 11273
rect -5240 11123 -5090 11273
rect -4880 11123 -4730 11273
rect -4520 11123 -4370 11273
rect -4160 11123 -4010 11273
rect -3800 11123 -3650 11273
rect -3440 11123 -3290 11273
rect -3080 11123 -2930 11273
rect -2720 11123 -2570 11273
rect -2360 11123 -2210 11273
rect -2000 11123 -1850 11273
rect -1640 11123 -1490 11273
rect -1280 11123 -1130 11273
rect -920 11123 -770 11273
rect -560 11123 -410 11273
rect -8840 10763 -8690 10913
rect -8480 10763 -8330 10913
rect -8120 10763 -7970 10913
rect -7760 10763 -7610 10913
rect -7400 10763 -7250 10913
rect -7040 10763 -6890 10913
rect -6680 10763 -6530 10913
rect -6320 10763 -6170 10913
rect -5960 10763 -5810 10913
rect -5600 10763 -5450 10913
rect -5240 10763 -5090 10913
rect -4880 10763 -4730 10913
rect -4520 10763 -4370 10913
rect -4160 10763 -4010 10913
rect -3800 10763 -3650 10913
rect -3440 10763 -3290 10913
rect -3080 10763 -2930 10913
rect -2720 10763 -2570 10913
rect -2360 10763 -2210 10913
rect -2000 10763 -1850 10913
rect -9560 11483 -9410 11633
rect -1640 10763 -1490 10913
rect -9200 11483 -9050 11633
rect -1280 10763 -1130 10913
rect -8840 11483 -8690 11633
rect -920 10763 -770 10913
rect -8480 11483 -8330 11633
rect -560 10763 -410 10913
rect -8120 11483 -7970 11633
rect -9560 10763 -9410 10913
rect -7760 11483 -7610 11633
rect -10280 10763 -10130 10913
rect -10280 11123 -10130 11273
rect -9920 10763 -9770 10913
rect -9920 11483 -9770 11633
rect -9920 11123 -9770 11273
rect -10280 11483 -10130 11633
rect -18560 11483 -18410 11633
rect -18920 10763 -18770 10913
rect -17120 11123 -16970 11273
rect -13520 11483 -13370 11633
rect -16760 11123 -16610 11273
rect -19280 11123 -19130 11273
rect -10640 10763 -10490 10913
rect -16400 11123 -16250 11273
rect -13160 11483 -13010 11633
rect -18560 10763 -18410 10913
rect -16040 11123 -15890 11273
rect -15320 10763 -15170 10913
rect -18200 11483 -18050 11633
rect -15680 11483 -15530 11633
rect -12800 10763 -12650 10913
rect -15680 11123 -15530 11273
rect -14600 10763 -14450 10913
rect -18200 10763 -18050 10913
rect -12800 11483 -12650 11633
rect -13520 10763 -13370 10913
rect -15320 11123 -15170 11273
rect -11720 10763 -11570 10913
rect -16760 11483 -16610 11633
rect -10640 11123 -10490 11273
rect -18920 11123 -18770 11273
rect -17840 10763 -17690 10913
rect -14960 11123 -14810 11273
rect -19640 11123 -19490 11273
rect -13880 11483 -13730 11633
rect -19640 11483 -19490 11633
rect -12440 11483 -12290 11633
rect -17120 11483 -16970 11633
rect -14600 11123 -14450 11273
rect -18200 11123 -18050 11273
rect -17840 11483 -17690 11633
rect -18560 11123 -18410 11273
rect -14240 11123 -14090 11273
rect -13160 10763 -13010 10913
rect -11000 11483 -10850 11633
rect -12080 11483 -11930 11633
rect -15320 11483 -15170 11633
rect -18920 11483 -18770 11633
rect -16400 11483 -16250 11633
rect -13880 11123 -13730 11273
rect -17480 10763 -17330 10913
rect -17480 11123 -17330 11273
rect -14240 10763 -14090 10913
rect -11360 11123 -11210 11273
rect -19280 11483 -19130 11633
rect -19640 10763 -19490 10913
rect -14960 10763 -14810 10913
rect -13520 11123 -13370 11273
rect -17120 10763 -16970 10913
rect -12080 11123 -11930 11273
rect -11000 10763 -10850 10913
rect -11720 11483 -11570 11633
rect -14960 11483 -14810 11633
rect -12080 10763 -11930 10913
rect -10640 11483 -10490 11633
rect -13160 11123 -13010 11273
rect -16760 10763 -16610 10913
rect -15680 10763 -15530 10913
rect -11720 11123 -11570 11273
rect -17480 11483 -17330 11633
rect -11360 10763 -11210 10913
rect -19280 10763 -19130 10913
rect -13880 10763 -13730 10913
rect -12800 11123 -12650 11273
rect -16400 10763 -16250 10913
rect -12440 10763 -12290 10913
rect -14240 11483 -14090 11633
rect -11360 11483 -11210 11633
rect -14600 11483 -14450 11633
rect -16040 11483 -15890 11633
rect -11000 11123 -10850 11273
rect -12440 11123 -12290 11273
rect -16040 10763 -15890 10913
rect -17840 11123 -17690 11273
rect -19235 -185 -19085 -35
rect -19605 -555 -19455 -405
rect -19235 -555 -19085 -405
rect -19605 -185 -19455 -35
<< l69d20 >>
rect -19690 -640 -19000 50
rect -19725 10678 20195 11718
<< l69d16 >>
rect -19690 -640 -19000 50
rect -19725 10678 20195 11718
<< labels >>
rlabel l68d5 -20211 188 -20211 188 0 CTRL
rlabel l68d5 19980 4475 19980 4475 0 OUT
rlabel l68d5 -19260 4545 -19260 4545 0 OUT
rlabel l68d5 890 4535 890 4535 0 OUT
rlabel l68d5 11225 4570 11225 4570 0 OUT
rlabel l68d5 -10320 4715 -10320 4715 0 OUT
rlabel l68d5 -20310 9300 -20310 9300 0 IN
rlabel l68d5 -20315 1665 -20315 1665 0 IN
rlabel l68d5 -20310 6100 -20310 6100 0 IN
rlabel l68d5 -20310 7935 -20310 7935 0 IN
rlabel l68d5 -20300 4170 -20300 4170 0 IN
rlabel l69d5 -19355 -235 -19355 -235 0 VSS
rlabel l69d5 -19365 11230 -19365 11230 0 VDD
rlabel l69d5 19970 11215 19970 11215 0 VDD
rlabel l69d5 45 11185 45 11185 0 VDD
rlabel l69d5 11760 11145 11760 11145 0 VDD
rlabel l69d5 -10080 11250 -10080 11250 0 VDD
use nfetx2410 nfetx2410_1
timestamp 1698899266
transform 0 -1 10235 1 0 745
box -125 -200 3445 30540
use pfetx246 pfetx246_1
timestamp 1698899266
transform 0 -1 20235 1 0 4495
box -305 -380 7671 40720
use nfet nfet_1
timestamp 1698899266
transform 0 -1 -18845 -1 0 585
box -125 -200 1374 1540
<< end >>
