magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< nwell >>
rect 0 0 1595 8220
<< pmos >>
rect 265 76 1065 8076
<< pdiff >>
rect 61 8053 265 8076
rect 61 8019 74 8053
rect 108 8019 146 8053
rect 180 8019 218 8053
rect 252 8019 265 8053
rect 61 7981 265 8019
rect 61 7947 74 7981
rect 108 7947 146 7981
rect 180 7947 218 7981
rect 252 7947 265 7981
rect 61 7909 265 7947
rect 61 7875 74 7909
rect 108 7875 146 7909
rect 180 7875 218 7909
rect 252 7875 265 7909
rect 61 7837 265 7875
rect 61 7803 74 7837
rect 108 7803 146 7837
rect 180 7803 218 7837
rect 252 7803 265 7837
rect 61 7765 265 7803
rect 61 7731 74 7765
rect 108 7731 146 7765
rect 180 7731 218 7765
rect 252 7731 265 7765
rect 61 7693 265 7731
rect 61 7659 74 7693
rect 108 7659 146 7693
rect 180 7659 218 7693
rect 252 7659 265 7693
rect 61 7621 265 7659
rect 61 7587 74 7621
rect 108 7587 146 7621
rect 180 7587 218 7621
rect 252 7587 265 7621
rect 61 7549 265 7587
rect 61 7515 74 7549
rect 108 7515 146 7549
rect 180 7515 218 7549
rect 252 7515 265 7549
rect 61 7477 265 7515
rect 61 7443 74 7477
rect 108 7443 146 7477
rect 180 7443 218 7477
rect 252 7443 265 7477
rect 61 7405 265 7443
rect 61 7371 74 7405
rect 108 7371 146 7405
rect 180 7371 218 7405
rect 252 7371 265 7405
rect 61 7333 265 7371
rect 61 7299 74 7333
rect 108 7299 146 7333
rect 180 7299 218 7333
rect 252 7299 265 7333
rect 61 7261 265 7299
rect 61 7227 74 7261
rect 108 7227 146 7261
rect 180 7227 218 7261
rect 252 7227 265 7261
rect 61 7189 265 7227
rect 61 7155 74 7189
rect 108 7155 146 7189
rect 180 7155 218 7189
rect 252 7155 265 7189
rect 61 7117 265 7155
rect 61 7083 74 7117
rect 108 7083 146 7117
rect 180 7083 218 7117
rect 252 7083 265 7117
rect 61 7045 265 7083
rect 61 7011 74 7045
rect 108 7011 146 7045
rect 180 7011 218 7045
rect 252 7011 265 7045
rect 61 6973 265 7011
rect 61 6939 74 6973
rect 108 6939 146 6973
rect 180 6939 218 6973
rect 252 6939 265 6973
rect 61 6901 265 6939
rect 61 6867 74 6901
rect 108 6867 146 6901
rect 180 6867 218 6901
rect 252 6867 265 6901
rect 61 6829 265 6867
rect 61 6795 74 6829
rect 108 6795 146 6829
rect 180 6795 218 6829
rect 252 6795 265 6829
rect 61 6757 265 6795
rect 61 6723 74 6757
rect 108 6723 146 6757
rect 180 6723 218 6757
rect 252 6723 265 6757
rect 61 6685 265 6723
rect 61 6651 74 6685
rect 108 6651 146 6685
rect 180 6651 218 6685
rect 252 6651 265 6685
rect 61 6613 265 6651
rect 61 6579 74 6613
rect 108 6579 146 6613
rect 180 6579 218 6613
rect 252 6579 265 6613
rect 61 6541 265 6579
rect 61 6507 74 6541
rect 108 6507 146 6541
rect 180 6507 218 6541
rect 252 6507 265 6541
rect 61 6469 265 6507
rect 61 6435 74 6469
rect 108 6435 146 6469
rect 180 6435 218 6469
rect 252 6435 265 6469
rect 61 6397 265 6435
rect 61 6363 74 6397
rect 108 6363 146 6397
rect 180 6363 218 6397
rect 252 6363 265 6397
rect 61 6325 265 6363
rect 61 6291 74 6325
rect 108 6291 146 6325
rect 180 6291 218 6325
rect 252 6291 265 6325
rect 61 6253 265 6291
rect 61 6219 74 6253
rect 108 6219 146 6253
rect 180 6219 218 6253
rect 252 6219 265 6253
rect 61 6181 265 6219
rect 61 6147 74 6181
rect 108 6147 146 6181
rect 180 6147 218 6181
rect 252 6147 265 6181
rect 61 6109 265 6147
rect 61 6075 74 6109
rect 108 6075 146 6109
rect 180 6075 218 6109
rect 252 6075 265 6109
rect 61 6037 265 6075
rect 61 6003 74 6037
rect 108 6003 146 6037
rect 180 6003 218 6037
rect 252 6003 265 6037
rect 61 5965 265 6003
rect 61 5931 74 5965
rect 108 5931 146 5965
rect 180 5931 218 5965
rect 252 5931 265 5965
rect 61 5893 265 5931
rect 61 5859 74 5893
rect 108 5859 146 5893
rect 180 5859 218 5893
rect 252 5859 265 5893
rect 61 5821 265 5859
rect 61 5787 74 5821
rect 108 5787 146 5821
rect 180 5787 218 5821
rect 252 5787 265 5821
rect 61 5749 265 5787
rect 61 5715 74 5749
rect 108 5715 146 5749
rect 180 5715 218 5749
rect 252 5715 265 5749
rect 61 5677 265 5715
rect 61 5643 74 5677
rect 108 5643 146 5677
rect 180 5643 218 5677
rect 252 5643 265 5677
rect 61 5605 265 5643
rect 61 5571 74 5605
rect 108 5571 146 5605
rect 180 5571 218 5605
rect 252 5571 265 5605
rect 61 5533 265 5571
rect 61 5499 74 5533
rect 108 5499 146 5533
rect 180 5499 218 5533
rect 252 5499 265 5533
rect 61 5461 265 5499
rect 61 5427 74 5461
rect 108 5427 146 5461
rect 180 5427 218 5461
rect 252 5427 265 5461
rect 61 5389 265 5427
rect 61 5355 74 5389
rect 108 5355 146 5389
rect 180 5355 218 5389
rect 252 5355 265 5389
rect 61 5317 265 5355
rect 61 5283 74 5317
rect 108 5283 146 5317
rect 180 5283 218 5317
rect 252 5283 265 5317
rect 61 5245 265 5283
rect 61 5211 74 5245
rect 108 5211 146 5245
rect 180 5211 218 5245
rect 252 5211 265 5245
rect 61 5173 265 5211
rect 61 5139 74 5173
rect 108 5139 146 5173
rect 180 5139 218 5173
rect 252 5139 265 5173
rect 61 5101 265 5139
rect 61 5067 74 5101
rect 108 5067 146 5101
rect 180 5067 218 5101
rect 252 5067 265 5101
rect 61 5029 265 5067
rect 61 4995 74 5029
rect 108 4995 146 5029
rect 180 4995 218 5029
rect 252 4995 265 5029
rect 61 4957 265 4995
rect 61 4923 74 4957
rect 108 4923 146 4957
rect 180 4923 218 4957
rect 252 4923 265 4957
rect 61 4885 265 4923
rect 61 4851 74 4885
rect 108 4851 146 4885
rect 180 4851 218 4885
rect 252 4851 265 4885
rect 61 4813 265 4851
rect 61 4779 74 4813
rect 108 4779 146 4813
rect 180 4779 218 4813
rect 252 4779 265 4813
rect 61 4741 265 4779
rect 61 4707 74 4741
rect 108 4707 146 4741
rect 180 4707 218 4741
rect 252 4707 265 4741
rect 61 4669 265 4707
rect 61 4635 74 4669
rect 108 4635 146 4669
rect 180 4635 218 4669
rect 252 4635 265 4669
rect 61 4597 265 4635
rect 61 4563 74 4597
rect 108 4563 146 4597
rect 180 4563 218 4597
rect 252 4563 265 4597
rect 61 4525 265 4563
rect 61 4491 74 4525
rect 108 4491 146 4525
rect 180 4491 218 4525
rect 252 4491 265 4525
rect 61 4453 265 4491
rect 61 4419 74 4453
rect 108 4419 146 4453
rect 180 4419 218 4453
rect 252 4419 265 4453
rect 61 4381 265 4419
rect 61 4347 74 4381
rect 108 4347 146 4381
rect 180 4347 218 4381
rect 252 4347 265 4381
rect 61 4309 265 4347
rect 61 4275 74 4309
rect 108 4275 146 4309
rect 180 4275 218 4309
rect 252 4275 265 4309
rect 61 4237 265 4275
rect 61 4203 74 4237
rect 108 4203 146 4237
rect 180 4203 218 4237
rect 252 4203 265 4237
rect 61 4165 265 4203
rect 61 4131 74 4165
rect 108 4131 146 4165
rect 180 4131 218 4165
rect 252 4131 265 4165
rect 61 4093 265 4131
rect 61 4059 74 4093
rect 108 4059 146 4093
rect 180 4059 218 4093
rect 252 4059 265 4093
rect 61 4021 265 4059
rect 61 3987 74 4021
rect 108 3987 146 4021
rect 180 3987 218 4021
rect 252 3987 265 4021
rect 61 3949 265 3987
rect 61 3915 74 3949
rect 108 3915 146 3949
rect 180 3915 218 3949
rect 252 3915 265 3949
rect 61 3877 265 3915
rect 61 3843 74 3877
rect 108 3843 146 3877
rect 180 3843 218 3877
rect 252 3843 265 3877
rect 61 3805 265 3843
rect 61 3771 74 3805
rect 108 3771 146 3805
rect 180 3771 218 3805
rect 252 3771 265 3805
rect 61 3733 265 3771
rect 61 3699 74 3733
rect 108 3699 146 3733
rect 180 3699 218 3733
rect 252 3699 265 3733
rect 61 3661 265 3699
rect 61 3627 74 3661
rect 108 3627 146 3661
rect 180 3627 218 3661
rect 252 3627 265 3661
rect 61 3589 265 3627
rect 61 3555 74 3589
rect 108 3555 146 3589
rect 180 3555 218 3589
rect 252 3555 265 3589
rect 61 3517 265 3555
rect 61 3483 74 3517
rect 108 3483 146 3517
rect 180 3483 218 3517
rect 252 3483 265 3517
rect 61 3445 265 3483
rect 61 3411 74 3445
rect 108 3411 146 3445
rect 180 3411 218 3445
rect 252 3411 265 3445
rect 61 3373 265 3411
rect 61 3339 74 3373
rect 108 3339 146 3373
rect 180 3339 218 3373
rect 252 3339 265 3373
rect 61 3301 265 3339
rect 61 3267 74 3301
rect 108 3267 146 3301
rect 180 3267 218 3301
rect 252 3267 265 3301
rect 61 3229 265 3267
rect 61 3195 74 3229
rect 108 3195 146 3229
rect 180 3195 218 3229
rect 252 3195 265 3229
rect 61 3157 265 3195
rect 61 3123 74 3157
rect 108 3123 146 3157
rect 180 3123 218 3157
rect 252 3123 265 3157
rect 61 3085 265 3123
rect 61 3051 74 3085
rect 108 3051 146 3085
rect 180 3051 218 3085
rect 252 3051 265 3085
rect 61 3013 265 3051
rect 61 2979 74 3013
rect 108 2979 146 3013
rect 180 2979 218 3013
rect 252 2979 265 3013
rect 61 2941 265 2979
rect 61 2907 74 2941
rect 108 2907 146 2941
rect 180 2907 218 2941
rect 252 2907 265 2941
rect 61 2869 265 2907
rect 61 2835 74 2869
rect 108 2835 146 2869
rect 180 2835 218 2869
rect 252 2835 265 2869
rect 61 2797 265 2835
rect 61 2763 74 2797
rect 108 2763 146 2797
rect 180 2763 218 2797
rect 252 2763 265 2797
rect 61 2725 265 2763
rect 61 2691 74 2725
rect 108 2691 146 2725
rect 180 2691 218 2725
rect 252 2691 265 2725
rect 61 2653 265 2691
rect 61 2619 74 2653
rect 108 2619 146 2653
rect 180 2619 218 2653
rect 252 2619 265 2653
rect 61 2581 265 2619
rect 61 2547 74 2581
rect 108 2547 146 2581
rect 180 2547 218 2581
rect 252 2547 265 2581
rect 61 2509 265 2547
rect 61 2475 74 2509
rect 108 2475 146 2509
rect 180 2475 218 2509
rect 252 2475 265 2509
rect 61 2437 265 2475
rect 61 2403 74 2437
rect 108 2403 146 2437
rect 180 2403 218 2437
rect 252 2403 265 2437
rect 61 2365 265 2403
rect 61 2331 74 2365
rect 108 2331 146 2365
rect 180 2331 218 2365
rect 252 2331 265 2365
rect 61 2293 265 2331
rect 61 2259 74 2293
rect 108 2259 146 2293
rect 180 2259 218 2293
rect 252 2259 265 2293
rect 61 2221 265 2259
rect 61 2187 74 2221
rect 108 2187 146 2221
rect 180 2187 218 2221
rect 252 2187 265 2221
rect 61 2149 265 2187
rect 61 2115 74 2149
rect 108 2115 146 2149
rect 180 2115 218 2149
rect 252 2115 265 2149
rect 61 2077 265 2115
rect 61 2043 74 2077
rect 108 2043 146 2077
rect 180 2043 218 2077
rect 252 2043 265 2077
rect 61 2005 265 2043
rect 61 1971 74 2005
rect 108 1971 146 2005
rect 180 1971 218 2005
rect 252 1971 265 2005
rect 61 1933 265 1971
rect 61 1899 74 1933
rect 108 1899 146 1933
rect 180 1899 218 1933
rect 252 1899 265 1933
rect 61 1861 265 1899
rect 61 1827 74 1861
rect 108 1827 146 1861
rect 180 1827 218 1861
rect 252 1827 265 1861
rect 61 1789 265 1827
rect 61 1755 74 1789
rect 108 1755 146 1789
rect 180 1755 218 1789
rect 252 1755 265 1789
rect 61 1717 265 1755
rect 61 1683 74 1717
rect 108 1683 146 1717
rect 180 1683 218 1717
rect 252 1683 265 1717
rect 61 1645 265 1683
rect 61 1611 74 1645
rect 108 1611 146 1645
rect 180 1611 218 1645
rect 252 1611 265 1645
rect 61 1573 265 1611
rect 61 1539 74 1573
rect 108 1539 146 1573
rect 180 1539 218 1573
rect 252 1539 265 1573
rect 61 1501 265 1539
rect 61 1467 74 1501
rect 108 1467 146 1501
rect 180 1467 218 1501
rect 252 1467 265 1501
rect 61 1429 265 1467
rect 61 1395 74 1429
rect 108 1395 146 1429
rect 180 1395 218 1429
rect 252 1395 265 1429
rect 61 1357 265 1395
rect 61 1323 74 1357
rect 108 1323 146 1357
rect 180 1323 218 1357
rect 252 1323 265 1357
rect 61 1285 265 1323
rect 61 1251 74 1285
rect 108 1251 146 1285
rect 180 1251 218 1285
rect 252 1251 265 1285
rect 61 1213 265 1251
rect 61 1179 74 1213
rect 108 1179 146 1213
rect 180 1179 218 1213
rect 252 1179 265 1213
rect 61 1141 265 1179
rect 61 1107 74 1141
rect 108 1107 146 1141
rect 180 1107 218 1141
rect 252 1107 265 1141
rect 61 1069 265 1107
rect 61 1035 74 1069
rect 108 1035 146 1069
rect 180 1035 218 1069
rect 252 1035 265 1069
rect 61 997 265 1035
rect 61 963 74 997
rect 108 963 146 997
rect 180 963 218 997
rect 252 963 265 997
rect 61 925 265 963
rect 61 891 74 925
rect 108 891 146 925
rect 180 891 218 925
rect 252 891 265 925
rect 61 853 265 891
rect 61 819 74 853
rect 108 819 146 853
rect 180 819 218 853
rect 252 819 265 853
rect 61 781 265 819
rect 61 747 74 781
rect 108 747 146 781
rect 180 747 218 781
rect 252 747 265 781
rect 61 709 265 747
rect 61 675 74 709
rect 108 675 146 709
rect 180 675 218 709
rect 252 675 265 709
rect 61 637 265 675
rect 61 603 74 637
rect 108 603 146 637
rect 180 603 218 637
rect 252 603 265 637
rect 61 565 265 603
rect 61 531 74 565
rect 108 531 146 565
rect 180 531 218 565
rect 252 531 265 565
rect 61 493 265 531
rect 61 459 74 493
rect 108 459 146 493
rect 180 459 218 493
rect 252 459 265 493
rect 61 421 265 459
rect 61 387 74 421
rect 108 387 146 421
rect 180 387 218 421
rect 252 387 265 421
rect 61 349 265 387
rect 61 315 74 349
rect 108 315 146 349
rect 180 315 218 349
rect 252 315 265 349
rect 61 277 265 315
rect 61 243 74 277
rect 108 243 146 277
rect 180 243 218 277
rect 252 243 265 277
rect 61 205 265 243
rect 61 171 74 205
rect 108 171 146 205
rect 180 171 218 205
rect 252 171 265 205
rect 61 133 265 171
rect 61 99 74 133
rect 108 99 146 133
rect 180 99 218 133
rect 252 99 265 133
rect 61 76 265 99
rect 1065 8053 1269 8076
rect 1065 8019 1078 8053
rect 1112 8019 1150 8053
rect 1184 8019 1222 8053
rect 1256 8019 1269 8053
rect 1065 7981 1269 8019
rect 1065 7947 1078 7981
rect 1112 7947 1150 7981
rect 1184 7947 1222 7981
rect 1256 7947 1269 7981
rect 1065 7909 1269 7947
rect 1065 7875 1078 7909
rect 1112 7875 1150 7909
rect 1184 7875 1222 7909
rect 1256 7875 1269 7909
rect 1065 7837 1269 7875
rect 1065 7803 1078 7837
rect 1112 7803 1150 7837
rect 1184 7803 1222 7837
rect 1256 7803 1269 7837
rect 1065 7765 1269 7803
rect 1065 7731 1078 7765
rect 1112 7731 1150 7765
rect 1184 7731 1222 7765
rect 1256 7731 1269 7765
rect 1065 7693 1269 7731
rect 1065 7659 1078 7693
rect 1112 7659 1150 7693
rect 1184 7659 1222 7693
rect 1256 7659 1269 7693
rect 1065 7621 1269 7659
rect 1065 7587 1078 7621
rect 1112 7587 1150 7621
rect 1184 7587 1222 7621
rect 1256 7587 1269 7621
rect 1065 7549 1269 7587
rect 1065 7515 1078 7549
rect 1112 7515 1150 7549
rect 1184 7515 1222 7549
rect 1256 7515 1269 7549
rect 1065 7477 1269 7515
rect 1065 7443 1078 7477
rect 1112 7443 1150 7477
rect 1184 7443 1222 7477
rect 1256 7443 1269 7477
rect 1065 7405 1269 7443
rect 1065 7371 1078 7405
rect 1112 7371 1150 7405
rect 1184 7371 1222 7405
rect 1256 7371 1269 7405
rect 1065 7333 1269 7371
rect 1065 7299 1078 7333
rect 1112 7299 1150 7333
rect 1184 7299 1222 7333
rect 1256 7299 1269 7333
rect 1065 7261 1269 7299
rect 1065 7227 1078 7261
rect 1112 7227 1150 7261
rect 1184 7227 1222 7261
rect 1256 7227 1269 7261
rect 1065 7189 1269 7227
rect 1065 7155 1078 7189
rect 1112 7155 1150 7189
rect 1184 7155 1222 7189
rect 1256 7155 1269 7189
rect 1065 7117 1269 7155
rect 1065 7083 1078 7117
rect 1112 7083 1150 7117
rect 1184 7083 1222 7117
rect 1256 7083 1269 7117
rect 1065 7045 1269 7083
rect 1065 7011 1078 7045
rect 1112 7011 1150 7045
rect 1184 7011 1222 7045
rect 1256 7011 1269 7045
rect 1065 6973 1269 7011
rect 1065 6939 1078 6973
rect 1112 6939 1150 6973
rect 1184 6939 1222 6973
rect 1256 6939 1269 6973
rect 1065 6901 1269 6939
rect 1065 6867 1078 6901
rect 1112 6867 1150 6901
rect 1184 6867 1222 6901
rect 1256 6867 1269 6901
rect 1065 6829 1269 6867
rect 1065 6795 1078 6829
rect 1112 6795 1150 6829
rect 1184 6795 1222 6829
rect 1256 6795 1269 6829
rect 1065 6757 1269 6795
rect 1065 6723 1078 6757
rect 1112 6723 1150 6757
rect 1184 6723 1222 6757
rect 1256 6723 1269 6757
rect 1065 6685 1269 6723
rect 1065 6651 1078 6685
rect 1112 6651 1150 6685
rect 1184 6651 1222 6685
rect 1256 6651 1269 6685
rect 1065 6613 1269 6651
rect 1065 6579 1078 6613
rect 1112 6579 1150 6613
rect 1184 6579 1222 6613
rect 1256 6579 1269 6613
rect 1065 6541 1269 6579
rect 1065 6507 1078 6541
rect 1112 6507 1150 6541
rect 1184 6507 1222 6541
rect 1256 6507 1269 6541
rect 1065 6469 1269 6507
rect 1065 6435 1078 6469
rect 1112 6435 1150 6469
rect 1184 6435 1222 6469
rect 1256 6435 1269 6469
rect 1065 6397 1269 6435
rect 1065 6363 1078 6397
rect 1112 6363 1150 6397
rect 1184 6363 1222 6397
rect 1256 6363 1269 6397
rect 1065 6325 1269 6363
rect 1065 6291 1078 6325
rect 1112 6291 1150 6325
rect 1184 6291 1222 6325
rect 1256 6291 1269 6325
rect 1065 6253 1269 6291
rect 1065 6219 1078 6253
rect 1112 6219 1150 6253
rect 1184 6219 1222 6253
rect 1256 6219 1269 6253
rect 1065 6181 1269 6219
rect 1065 6147 1078 6181
rect 1112 6147 1150 6181
rect 1184 6147 1222 6181
rect 1256 6147 1269 6181
rect 1065 6109 1269 6147
rect 1065 6075 1078 6109
rect 1112 6075 1150 6109
rect 1184 6075 1222 6109
rect 1256 6075 1269 6109
rect 1065 6037 1269 6075
rect 1065 6003 1078 6037
rect 1112 6003 1150 6037
rect 1184 6003 1222 6037
rect 1256 6003 1269 6037
rect 1065 5965 1269 6003
rect 1065 5931 1078 5965
rect 1112 5931 1150 5965
rect 1184 5931 1222 5965
rect 1256 5931 1269 5965
rect 1065 5893 1269 5931
rect 1065 5859 1078 5893
rect 1112 5859 1150 5893
rect 1184 5859 1222 5893
rect 1256 5859 1269 5893
rect 1065 5821 1269 5859
rect 1065 5787 1078 5821
rect 1112 5787 1150 5821
rect 1184 5787 1222 5821
rect 1256 5787 1269 5821
rect 1065 5749 1269 5787
rect 1065 5715 1078 5749
rect 1112 5715 1150 5749
rect 1184 5715 1222 5749
rect 1256 5715 1269 5749
rect 1065 5677 1269 5715
rect 1065 5643 1078 5677
rect 1112 5643 1150 5677
rect 1184 5643 1222 5677
rect 1256 5643 1269 5677
rect 1065 5605 1269 5643
rect 1065 5571 1078 5605
rect 1112 5571 1150 5605
rect 1184 5571 1222 5605
rect 1256 5571 1269 5605
rect 1065 5533 1269 5571
rect 1065 5499 1078 5533
rect 1112 5499 1150 5533
rect 1184 5499 1222 5533
rect 1256 5499 1269 5533
rect 1065 5461 1269 5499
rect 1065 5427 1078 5461
rect 1112 5427 1150 5461
rect 1184 5427 1222 5461
rect 1256 5427 1269 5461
rect 1065 5389 1269 5427
rect 1065 5355 1078 5389
rect 1112 5355 1150 5389
rect 1184 5355 1222 5389
rect 1256 5355 1269 5389
rect 1065 5317 1269 5355
rect 1065 5283 1078 5317
rect 1112 5283 1150 5317
rect 1184 5283 1222 5317
rect 1256 5283 1269 5317
rect 1065 5245 1269 5283
rect 1065 5211 1078 5245
rect 1112 5211 1150 5245
rect 1184 5211 1222 5245
rect 1256 5211 1269 5245
rect 1065 5173 1269 5211
rect 1065 5139 1078 5173
rect 1112 5139 1150 5173
rect 1184 5139 1222 5173
rect 1256 5139 1269 5173
rect 1065 5101 1269 5139
rect 1065 5067 1078 5101
rect 1112 5067 1150 5101
rect 1184 5067 1222 5101
rect 1256 5067 1269 5101
rect 1065 5029 1269 5067
rect 1065 4995 1078 5029
rect 1112 4995 1150 5029
rect 1184 4995 1222 5029
rect 1256 4995 1269 5029
rect 1065 4957 1269 4995
rect 1065 4923 1078 4957
rect 1112 4923 1150 4957
rect 1184 4923 1222 4957
rect 1256 4923 1269 4957
rect 1065 4885 1269 4923
rect 1065 4851 1078 4885
rect 1112 4851 1150 4885
rect 1184 4851 1222 4885
rect 1256 4851 1269 4885
rect 1065 4813 1269 4851
rect 1065 4779 1078 4813
rect 1112 4779 1150 4813
rect 1184 4779 1222 4813
rect 1256 4779 1269 4813
rect 1065 4741 1269 4779
rect 1065 4707 1078 4741
rect 1112 4707 1150 4741
rect 1184 4707 1222 4741
rect 1256 4707 1269 4741
rect 1065 4669 1269 4707
rect 1065 4635 1078 4669
rect 1112 4635 1150 4669
rect 1184 4635 1222 4669
rect 1256 4635 1269 4669
rect 1065 4597 1269 4635
rect 1065 4563 1078 4597
rect 1112 4563 1150 4597
rect 1184 4563 1222 4597
rect 1256 4563 1269 4597
rect 1065 4525 1269 4563
rect 1065 4491 1078 4525
rect 1112 4491 1150 4525
rect 1184 4491 1222 4525
rect 1256 4491 1269 4525
rect 1065 4453 1269 4491
rect 1065 4419 1078 4453
rect 1112 4419 1150 4453
rect 1184 4419 1222 4453
rect 1256 4419 1269 4453
rect 1065 4381 1269 4419
rect 1065 4347 1078 4381
rect 1112 4347 1150 4381
rect 1184 4347 1222 4381
rect 1256 4347 1269 4381
rect 1065 4309 1269 4347
rect 1065 4275 1078 4309
rect 1112 4275 1150 4309
rect 1184 4275 1222 4309
rect 1256 4275 1269 4309
rect 1065 4237 1269 4275
rect 1065 4203 1078 4237
rect 1112 4203 1150 4237
rect 1184 4203 1222 4237
rect 1256 4203 1269 4237
rect 1065 4165 1269 4203
rect 1065 4131 1078 4165
rect 1112 4131 1150 4165
rect 1184 4131 1222 4165
rect 1256 4131 1269 4165
rect 1065 4093 1269 4131
rect 1065 4059 1078 4093
rect 1112 4059 1150 4093
rect 1184 4059 1222 4093
rect 1256 4059 1269 4093
rect 1065 4021 1269 4059
rect 1065 3987 1078 4021
rect 1112 3987 1150 4021
rect 1184 3987 1222 4021
rect 1256 3987 1269 4021
rect 1065 3949 1269 3987
rect 1065 3915 1078 3949
rect 1112 3915 1150 3949
rect 1184 3915 1222 3949
rect 1256 3915 1269 3949
rect 1065 3877 1269 3915
rect 1065 3843 1078 3877
rect 1112 3843 1150 3877
rect 1184 3843 1222 3877
rect 1256 3843 1269 3877
rect 1065 3805 1269 3843
rect 1065 3771 1078 3805
rect 1112 3771 1150 3805
rect 1184 3771 1222 3805
rect 1256 3771 1269 3805
rect 1065 3733 1269 3771
rect 1065 3699 1078 3733
rect 1112 3699 1150 3733
rect 1184 3699 1222 3733
rect 1256 3699 1269 3733
rect 1065 3661 1269 3699
rect 1065 3627 1078 3661
rect 1112 3627 1150 3661
rect 1184 3627 1222 3661
rect 1256 3627 1269 3661
rect 1065 3589 1269 3627
rect 1065 3555 1078 3589
rect 1112 3555 1150 3589
rect 1184 3555 1222 3589
rect 1256 3555 1269 3589
rect 1065 3517 1269 3555
rect 1065 3483 1078 3517
rect 1112 3483 1150 3517
rect 1184 3483 1222 3517
rect 1256 3483 1269 3517
rect 1065 3445 1269 3483
rect 1065 3411 1078 3445
rect 1112 3411 1150 3445
rect 1184 3411 1222 3445
rect 1256 3411 1269 3445
rect 1065 3373 1269 3411
rect 1065 3339 1078 3373
rect 1112 3339 1150 3373
rect 1184 3339 1222 3373
rect 1256 3339 1269 3373
rect 1065 3301 1269 3339
rect 1065 3267 1078 3301
rect 1112 3267 1150 3301
rect 1184 3267 1222 3301
rect 1256 3267 1269 3301
rect 1065 3229 1269 3267
rect 1065 3195 1078 3229
rect 1112 3195 1150 3229
rect 1184 3195 1222 3229
rect 1256 3195 1269 3229
rect 1065 3157 1269 3195
rect 1065 3123 1078 3157
rect 1112 3123 1150 3157
rect 1184 3123 1222 3157
rect 1256 3123 1269 3157
rect 1065 3085 1269 3123
rect 1065 3051 1078 3085
rect 1112 3051 1150 3085
rect 1184 3051 1222 3085
rect 1256 3051 1269 3085
rect 1065 3013 1269 3051
rect 1065 2979 1078 3013
rect 1112 2979 1150 3013
rect 1184 2979 1222 3013
rect 1256 2979 1269 3013
rect 1065 2941 1269 2979
rect 1065 2907 1078 2941
rect 1112 2907 1150 2941
rect 1184 2907 1222 2941
rect 1256 2907 1269 2941
rect 1065 2869 1269 2907
rect 1065 2835 1078 2869
rect 1112 2835 1150 2869
rect 1184 2835 1222 2869
rect 1256 2835 1269 2869
rect 1065 2797 1269 2835
rect 1065 2763 1078 2797
rect 1112 2763 1150 2797
rect 1184 2763 1222 2797
rect 1256 2763 1269 2797
rect 1065 2725 1269 2763
rect 1065 2691 1078 2725
rect 1112 2691 1150 2725
rect 1184 2691 1222 2725
rect 1256 2691 1269 2725
rect 1065 2653 1269 2691
rect 1065 2619 1078 2653
rect 1112 2619 1150 2653
rect 1184 2619 1222 2653
rect 1256 2619 1269 2653
rect 1065 2581 1269 2619
rect 1065 2547 1078 2581
rect 1112 2547 1150 2581
rect 1184 2547 1222 2581
rect 1256 2547 1269 2581
rect 1065 2509 1269 2547
rect 1065 2475 1078 2509
rect 1112 2475 1150 2509
rect 1184 2475 1222 2509
rect 1256 2475 1269 2509
rect 1065 2437 1269 2475
rect 1065 2403 1078 2437
rect 1112 2403 1150 2437
rect 1184 2403 1222 2437
rect 1256 2403 1269 2437
rect 1065 2365 1269 2403
rect 1065 2331 1078 2365
rect 1112 2331 1150 2365
rect 1184 2331 1222 2365
rect 1256 2331 1269 2365
rect 1065 2293 1269 2331
rect 1065 2259 1078 2293
rect 1112 2259 1150 2293
rect 1184 2259 1222 2293
rect 1256 2259 1269 2293
rect 1065 2221 1269 2259
rect 1065 2187 1078 2221
rect 1112 2187 1150 2221
rect 1184 2187 1222 2221
rect 1256 2187 1269 2221
rect 1065 2149 1269 2187
rect 1065 2115 1078 2149
rect 1112 2115 1150 2149
rect 1184 2115 1222 2149
rect 1256 2115 1269 2149
rect 1065 2077 1269 2115
rect 1065 2043 1078 2077
rect 1112 2043 1150 2077
rect 1184 2043 1222 2077
rect 1256 2043 1269 2077
rect 1065 2005 1269 2043
rect 1065 1971 1078 2005
rect 1112 1971 1150 2005
rect 1184 1971 1222 2005
rect 1256 1971 1269 2005
rect 1065 1933 1269 1971
rect 1065 1899 1078 1933
rect 1112 1899 1150 1933
rect 1184 1899 1222 1933
rect 1256 1899 1269 1933
rect 1065 1861 1269 1899
rect 1065 1827 1078 1861
rect 1112 1827 1150 1861
rect 1184 1827 1222 1861
rect 1256 1827 1269 1861
rect 1065 1789 1269 1827
rect 1065 1755 1078 1789
rect 1112 1755 1150 1789
rect 1184 1755 1222 1789
rect 1256 1755 1269 1789
rect 1065 1717 1269 1755
rect 1065 1683 1078 1717
rect 1112 1683 1150 1717
rect 1184 1683 1222 1717
rect 1256 1683 1269 1717
rect 1065 1645 1269 1683
rect 1065 1611 1078 1645
rect 1112 1611 1150 1645
rect 1184 1611 1222 1645
rect 1256 1611 1269 1645
rect 1065 1573 1269 1611
rect 1065 1539 1078 1573
rect 1112 1539 1150 1573
rect 1184 1539 1222 1573
rect 1256 1539 1269 1573
rect 1065 1501 1269 1539
rect 1065 1467 1078 1501
rect 1112 1467 1150 1501
rect 1184 1467 1222 1501
rect 1256 1467 1269 1501
rect 1065 1429 1269 1467
rect 1065 1395 1078 1429
rect 1112 1395 1150 1429
rect 1184 1395 1222 1429
rect 1256 1395 1269 1429
rect 1065 1357 1269 1395
rect 1065 1323 1078 1357
rect 1112 1323 1150 1357
rect 1184 1323 1222 1357
rect 1256 1323 1269 1357
rect 1065 1285 1269 1323
rect 1065 1251 1078 1285
rect 1112 1251 1150 1285
rect 1184 1251 1222 1285
rect 1256 1251 1269 1285
rect 1065 1213 1269 1251
rect 1065 1179 1078 1213
rect 1112 1179 1150 1213
rect 1184 1179 1222 1213
rect 1256 1179 1269 1213
rect 1065 1141 1269 1179
rect 1065 1107 1078 1141
rect 1112 1107 1150 1141
rect 1184 1107 1222 1141
rect 1256 1107 1269 1141
rect 1065 1069 1269 1107
rect 1065 1035 1078 1069
rect 1112 1035 1150 1069
rect 1184 1035 1222 1069
rect 1256 1035 1269 1069
rect 1065 997 1269 1035
rect 1065 963 1078 997
rect 1112 963 1150 997
rect 1184 963 1222 997
rect 1256 963 1269 997
rect 1065 925 1269 963
rect 1065 891 1078 925
rect 1112 891 1150 925
rect 1184 891 1222 925
rect 1256 891 1269 925
rect 1065 853 1269 891
rect 1065 819 1078 853
rect 1112 819 1150 853
rect 1184 819 1222 853
rect 1256 819 1269 853
rect 1065 781 1269 819
rect 1065 747 1078 781
rect 1112 747 1150 781
rect 1184 747 1222 781
rect 1256 747 1269 781
rect 1065 709 1269 747
rect 1065 675 1078 709
rect 1112 675 1150 709
rect 1184 675 1222 709
rect 1256 675 1269 709
rect 1065 637 1269 675
rect 1065 603 1078 637
rect 1112 603 1150 637
rect 1184 603 1222 637
rect 1256 603 1269 637
rect 1065 565 1269 603
rect 1065 531 1078 565
rect 1112 531 1150 565
rect 1184 531 1222 565
rect 1256 531 1269 565
rect 1065 493 1269 531
rect 1065 459 1078 493
rect 1112 459 1150 493
rect 1184 459 1222 493
rect 1256 459 1269 493
rect 1065 421 1269 459
rect 1065 387 1078 421
rect 1112 387 1150 421
rect 1184 387 1222 421
rect 1256 387 1269 421
rect 1065 349 1269 387
rect 1065 315 1078 349
rect 1112 315 1150 349
rect 1184 315 1222 349
rect 1256 315 1269 349
rect 1065 277 1269 315
rect 1065 243 1078 277
rect 1112 243 1150 277
rect 1184 243 1222 277
rect 1256 243 1269 277
rect 1065 205 1269 243
rect 1065 171 1078 205
rect 1112 171 1150 205
rect 1184 171 1222 205
rect 1256 171 1269 205
rect 1065 133 1269 171
rect 1065 99 1078 133
rect 1112 99 1150 133
rect 1184 99 1222 133
rect 1256 99 1269 133
rect 1065 76 1269 99
<< pdiffc >>
rect 74 8019 108 8053
rect 146 8019 180 8053
rect 218 8019 252 8053
rect 74 7947 108 7981
rect 146 7947 180 7981
rect 218 7947 252 7981
rect 74 7875 108 7909
rect 146 7875 180 7909
rect 218 7875 252 7909
rect 74 7803 108 7837
rect 146 7803 180 7837
rect 218 7803 252 7837
rect 74 7731 108 7765
rect 146 7731 180 7765
rect 218 7731 252 7765
rect 74 7659 108 7693
rect 146 7659 180 7693
rect 218 7659 252 7693
rect 74 7587 108 7621
rect 146 7587 180 7621
rect 218 7587 252 7621
rect 74 7515 108 7549
rect 146 7515 180 7549
rect 218 7515 252 7549
rect 74 7443 108 7477
rect 146 7443 180 7477
rect 218 7443 252 7477
rect 74 7371 108 7405
rect 146 7371 180 7405
rect 218 7371 252 7405
rect 74 7299 108 7333
rect 146 7299 180 7333
rect 218 7299 252 7333
rect 74 7227 108 7261
rect 146 7227 180 7261
rect 218 7227 252 7261
rect 74 7155 108 7189
rect 146 7155 180 7189
rect 218 7155 252 7189
rect 74 7083 108 7117
rect 146 7083 180 7117
rect 218 7083 252 7117
rect 74 7011 108 7045
rect 146 7011 180 7045
rect 218 7011 252 7045
rect 74 6939 108 6973
rect 146 6939 180 6973
rect 218 6939 252 6973
rect 74 6867 108 6901
rect 146 6867 180 6901
rect 218 6867 252 6901
rect 74 6795 108 6829
rect 146 6795 180 6829
rect 218 6795 252 6829
rect 74 6723 108 6757
rect 146 6723 180 6757
rect 218 6723 252 6757
rect 74 6651 108 6685
rect 146 6651 180 6685
rect 218 6651 252 6685
rect 74 6579 108 6613
rect 146 6579 180 6613
rect 218 6579 252 6613
rect 74 6507 108 6541
rect 146 6507 180 6541
rect 218 6507 252 6541
rect 74 6435 108 6469
rect 146 6435 180 6469
rect 218 6435 252 6469
rect 74 6363 108 6397
rect 146 6363 180 6397
rect 218 6363 252 6397
rect 74 6291 108 6325
rect 146 6291 180 6325
rect 218 6291 252 6325
rect 74 6219 108 6253
rect 146 6219 180 6253
rect 218 6219 252 6253
rect 74 6147 108 6181
rect 146 6147 180 6181
rect 218 6147 252 6181
rect 74 6075 108 6109
rect 146 6075 180 6109
rect 218 6075 252 6109
rect 74 6003 108 6037
rect 146 6003 180 6037
rect 218 6003 252 6037
rect 74 5931 108 5965
rect 146 5931 180 5965
rect 218 5931 252 5965
rect 74 5859 108 5893
rect 146 5859 180 5893
rect 218 5859 252 5893
rect 74 5787 108 5821
rect 146 5787 180 5821
rect 218 5787 252 5821
rect 74 5715 108 5749
rect 146 5715 180 5749
rect 218 5715 252 5749
rect 74 5643 108 5677
rect 146 5643 180 5677
rect 218 5643 252 5677
rect 74 5571 108 5605
rect 146 5571 180 5605
rect 218 5571 252 5605
rect 74 5499 108 5533
rect 146 5499 180 5533
rect 218 5499 252 5533
rect 74 5427 108 5461
rect 146 5427 180 5461
rect 218 5427 252 5461
rect 74 5355 108 5389
rect 146 5355 180 5389
rect 218 5355 252 5389
rect 74 5283 108 5317
rect 146 5283 180 5317
rect 218 5283 252 5317
rect 74 5211 108 5245
rect 146 5211 180 5245
rect 218 5211 252 5245
rect 74 5139 108 5173
rect 146 5139 180 5173
rect 218 5139 252 5173
rect 74 5067 108 5101
rect 146 5067 180 5101
rect 218 5067 252 5101
rect 74 4995 108 5029
rect 146 4995 180 5029
rect 218 4995 252 5029
rect 74 4923 108 4957
rect 146 4923 180 4957
rect 218 4923 252 4957
rect 74 4851 108 4885
rect 146 4851 180 4885
rect 218 4851 252 4885
rect 74 4779 108 4813
rect 146 4779 180 4813
rect 218 4779 252 4813
rect 74 4707 108 4741
rect 146 4707 180 4741
rect 218 4707 252 4741
rect 74 4635 108 4669
rect 146 4635 180 4669
rect 218 4635 252 4669
rect 74 4563 108 4597
rect 146 4563 180 4597
rect 218 4563 252 4597
rect 74 4491 108 4525
rect 146 4491 180 4525
rect 218 4491 252 4525
rect 74 4419 108 4453
rect 146 4419 180 4453
rect 218 4419 252 4453
rect 74 4347 108 4381
rect 146 4347 180 4381
rect 218 4347 252 4381
rect 74 4275 108 4309
rect 146 4275 180 4309
rect 218 4275 252 4309
rect 74 4203 108 4237
rect 146 4203 180 4237
rect 218 4203 252 4237
rect 74 4131 108 4165
rect 146 4131 180 4165
rect 218 4131 252 4165
rect 74 4059 108 4093
rect 146 4059 180 4093
rect 218 4059 252 4093
rect 74 3987 108 4021
rect 146 3987 180 4021
rect 218 3987 252 4021
rect 74 3915 108 3949
rect 146 3915 180 3949
rect 218 3915 252 3949
rect 74 3843 108 3877
rect 146 3843 180 3877
rect 218 3843 252 3877
rect 74 3771 108 3805
rect 146 3771 180 3805
rect 218 3771 252 3805
rect 74 3699 108 3733
rect 146 3699 180 3733
rect 218 3699 252 3733
rect 74 3627 108 3661
rect 146 3627 180 3661
rect 218 3627 252 3661
rect 74 3555 108 3589
rect 146 3555 180 3589
rect 218 3555 252 3589
rect 74 3483 108 3517
rect 146 3483 180 3517
rect 218 3483 252 3517
rect 74 3411 108 3445
rect 146 3411 180 3445
rect 218 3411 252 3445
rect 74 3339 108 3373
rect 146 3339 180 3373
rect 218 3339 252 3373
rect 74 3267 108 3301
rect 146 3267 180 3301
rect 218 3267 252 3301
rect 74 3195 108 3229
rect 146 3195 180 3229
rect 218 3195 252 3229
rect 74 3123 108 3157
rect 146 3123 180 3157
rect 218 3123 252 3157
rect 74 3051 108 3085
rect 146 3051 180 3085
rect 218 3051 252 3085
rect 74 2979 108 3013
rect 146 2979 180 3013
rect 218 2979 252 3013
rect 74 2907 108 2941
rect 146 2907 180 2941
rect 218 2907 252 2941
rect 74 2835 108 2869
rect 146 2835 180 2869
rect 218 2835 252 2869
rect 74 2763 108 2797
rect 146 2763 180 2797
rect 218 2763 252 2797
rect 74 2691 108 2725
rect 146 2691 180 2725
rect 218 2691 252 2725
rect 74 2619 108 2653
rect 146 2619 180 2653
rect 218 2619 252 2653
rect 74 2547 108 2581
rect 146 2547 180 2581
rect 218 2547 252 2581
rect 74 2475 108 2509
rect 146 2475 180 2509
rect 218 2475 252 2509
rect 74 2403 108 2437
rect 146 2403 180 2437
rect 218 2403 252 2437
rect 74 2331 108 2365
rect 146 2331 180 2365
rect 218 2331 252 2365
rect 74 2259 108 2293
rect 146 2259 180 2293
rect 218 2259 252 2293
rect 74 2187 108 2221
rect 146 2187 180 2221
rect 218 2187 252 2221
rect 74 2115 108 2149
rect 146 2115 180 2149
rect 218 2115 252 2149
rect 74 2043 108 2077
rect 146 2043 180 2077
rect 218 2043 252 2077
rect 74 1971 108 2005
rect 146 1971 180 2005
rect 218 1971 252 2005
rect 74 1899 108 1933
rect 146 1899 180 1933
rect 218 1899 252 1933
rect 74 1827 108 1861
rect 146 1827 180 1861
rect 218 1827 252 1861
rect 74 1755 108 1789
rect 146 1755 180 1789
rect 218 1755 252 1789
rect 74 1683 108 1717
rect 146 1683 180 1717
rect 218 1683 252 1717
rect 74 1611 108 1645
rect 146 1611 180 1645
rect 218 1611 252 1645
rect 74 1539 108 1573
rect 146 1539 180 1573
rect 218 1539 252 1573
rect 74 1467 108 1501
rect 146 1467 180 1501
rect 218 1467 252 1501
rect 74 1395 108 1429
rect 146 1395 180 1429
rect 218 1395 252 1429
rect 74 1323 108 1357
rect 146 1323 180 1357
rect 218 1323 252 1357
rect 74 1251 108 1285
rect 146 1251 180 1285
rect 218 1251 252 1285
rect 74 1179 108 1213
rect 146 1179 180 1213
rect 218 1179 252 1213
rect 74 1107 108 1141
rect 146 1107 180 1141
rect 218 1107 252 1141
rect 74 1035 108 1069
rect 146 1035 180 1069
rect 218 1035 252 1069
rect 74 963 108 997
rect 146 963 180 997
rect 218 963 252 997
rect 74 891 108 925
rect 146 891 180 925
rect 218 891 252 925
rect 74 819 108 853
rect 146 819 180 853
rect 218 819 252 853
rect 74 747 108 781
rect 146 747 180 781
rect 218 747 252 781
rect 74 675 108 709
rect 146 675 180 709
rect 218 675 252 709
rect 74 603 108 637
rect 146 603 180 637
rect 218 603 252 637
rect 74 531 108 565
rect 146 531 180 565
rect 218 531 252 565
rect 74 459 108 493
rect 146 459 180 493
rect 218 459 252 493
rect 74 387 108 421
rect 146 387 180 421
rect 218 387 252 421
rect 74 315 108 349
rect 146 315 180 349
rect 218 315 252 349
rect 74 243 108 277
rect 146 243 180 277
rect 218 243 252 277
rect 74 171 108 205
rect 146 171 180 205
rect 218 171 252 205
rect 74 99 108 133
rect 146 99 180 133
rect 218 99 252 133
rect 1078 8019 1112 8053
rect 1150 8019 1184 8053
rect 1222 8019 1256 8053
rect 1078 7947 1112 7981
rect 1150 7947 1184 7981
rect 1222 7947 1256 7981
rect 1078 7875 1112 7909
rect 1150 7875 1184 7909
rect 1222 7875 1256 7909
rect 1078 7803 1112 7837
rect 1150 7803 1184 7837
rect 1222 7803 1256 7837
rect 1078 7731 1112 7765
rect 1150 7731 1184 7765
rect 1222 7731 1256 7765
rect 1078 7659 1112 7693
rect 1150 7659 1184 7693
rect 1222 7659 1256 7693
rect 1078 7587 1112 7621
rect 1150 7587 1184 7621
rect 1222 7587 1256 7621
rect 1078 7515 1112 7549
rect 1150 7515 1184 7549
rect 1222 7515 1256 7549
rect 1078 7443 1112 7477
rect 1150 7443 1184 7477
rect 1222 7443 1256 7477
rect 1078 7371 1112 7405
rect 1150 7371 1184 7405
rect 1222 7371 1256 7405
rect 1078 7299 1112 7333
rect 1150 7299 1184 7333
rect 1222 7299 1256 7333
rect 1078 7227 1112 7261
rect 1150 7227 1184 7261
rect 1222 7227 1256 7261
rect 1078 7155 1112 7189
rect 1150 7155 1184 7189
rect 1222 7155 1256 7189
rect 1078 7083 1112 7117
rect 1150 7083 1184 7117
rect 1222 7083 1256 7117
rect 1078 7011 1112 7045
rect 1150 7011 1184 7045
rect 1222 7011 1256 7045
rect 1078 6939 1112 6973
rect 1150 6939 1184 6973
rect 1222 6939 1256 6973
rect 1078 6867 1112 6901
rect 1150 6867 1184 6901
rect 1222 6867 1256 6901
rect 1078 6795 1112 6829
rect 1150 6795 1184 6829
rect 1222 6795 1256 6829
rect 1078 6723 1112 6757
rect 1150 6723 1184 6757
rect 1222 6723 1256 6757
rect 1078 6651 1112 6685
rect 1150 6651 1184 6685
rect 1222 6651 1256 6685
rect 1078 6579 1112 6613
rect 1150 6579 1184 6613
rect 1222 6579 1256 6613
rect 1078 6507 1112 6541
rect 1150 6507 1184 6541
rect 1222 6507 1256 6541
rect 1078 6435 1112 6469
rect 1150 6435 1184 6469
rect 1222 6435 1256 6469
rect 1078 6363 1112 6397
rect 1150 6363 1184 6397
rect 1222 6363 1256 6397
rect 1078 6291 1112 6325
rect 1150 6291 1184 6325
rect 1222 6291 1256 6325
rect 1078 6219 1112 6253
rect 1150 6219 1184 6253
rect 1222 6219 1256 6253
rect 1078 6147 1112 6181
rect 1150 6147 1184 6181
rect 1222 6147 1256 6181
rect 1078 6075 1112 6109
rect 1150 6075 1184 6109
rect 1222 6075 1256 6109
rect 1078 6003 1112 6037
rect 1150 6003 1184 6037
rect 1222 6003 1256 6037
rect 1078 5931 1112 5965
rect 1150 5931 1184 5965
rect 1222 5931 1256 5965
rect 1078 5859 1112 5893
rect 1150 5859 1184 5893
rect 1222 5859 1256 5893
rect 1078 5787 1112 5821
rect 1150 5787 1184 5821
rect 1222 5787 1256 5821
rect 1078 5715 1112 5749
rect 1150 5715 1184 5749
rect 1222 5715 1256 5749
rect 1078 5643 1112 5677
rect 1150 5643 1184 5677
rect 1222 5643 1256 5677
rect 1078 5571 1112 5605
rect 1150 5571 1184 5605
rect 1222 5571 1256 5605
rect 1078 5499 1112 5533
rect 1150 5499 1184 5533
rect 1222 5499 1256 5533
rect 1078 5427 1112 5461
rect 1150 5427 1184 5461
rect 1222 5427 1256 5461
rect 1078 5355 1112 5389
rect 1150 5355 1184 5389
rect 1222 5355 1256 5389
rect 1078 5283 1112 5317
rect 1150 5283 1184 5317
rect 1222 5283 1256 5317
rect 1078 5211 1112 5245
rect 1150 5211 1184 5245
rect 1222 5211 1256 5245
rect 1078 5139 1112 5173
rect 1150 5139 1184 5173
rect 1222 5139 1256 5173
rect 1078 5067 1112 5101
rect 1150 5067 1184 5101
rect 1222 5067 1256 5101
rect 1078 4995 1112 5029
rect 1150 4995 1184 5029
rect 1222 4995 1256 5029
rect 1078 4923 1112 4957
rect 1150 4923 1184 4957
rect 1222 4923 1256 4957
rect 1078 4851 1112 4885
rect 1150 4851 1184 4885
rect 1222 4851 1256 4885
rect 1078 4779 1112 4813
rect 1150 4779 1184 4813
rect 1222 4779 1256 4813
rect 1078 4707 1112 4741
rect 1150 4707 1184 4741
rect 1222 4707 1256 4741
rect 1078 4635 1112 4669
rect 1150 4635 1184 4669
rect 1222 4635 1256 4669
rect 1078 4563 1112 4597
rect 1150 4563 1184 4597
rect 1222 4563 1256 4597
rect 1078 4491 1112 4525
rect 1150 4491 1184 4525
rect 1222 4491 1256 4525
rect 1078 4419 1112 4453
rect 1150 4419 1184 4453
rect 1222 4419 1256 4453
rect 1078 4347 1112 4381
rect 1150 4347 1184 4381
rect 1222 4347 1256 4381
rect 1078 4275 1112 4309
rect 1150 4275 1184 4309
rect 1222 4275 1256 4309
rect 1078 4203 1112 4237
rect 1150 4203 1184 4237
rect 1222 4203 1256 4237
rect 1078 4131 1112 4165
rect 1150 4131 1184 4165
rect 1222 4131 1256 4165
rect 1078 4059 1112 4093
rect 1150 4059 1184 4093
rect 1222 4059 1256 4093
rect 1078 3987 1112 4021
rect 1150 3987 1184 4021
rect 1222 3987 1256 4021
rect 1078 3915 1112 3949
rect 1150 3915 1184 3949
rect 1222 3915 1256 3949
rect 1078 3843 1112 3877
rect 1150 3843 1184 3877
rect 1222 3843 1256 3877
rect 1078 3771 1112 3805
rect 1150 3771 1184 3805
rect 1222 3771 1256 3805
rect 1078 3699 1112 3733
rect 1150 3699 1184 3733
rect 1222 3699 1256 3733
rect 1078 3627 1112 3661
rect 1150 3627 1184 3661
rect 1222 3627 1256 3661
rect 1078 3555 1112 3589
rect 1150 3555 1184 3589
rect 1222 3555 1256 3589
rect 1078 3483 1112 3517
rect 1150 3483 1184 3517
rect 1222 3483 1256 3517
rect 1078 3411 1112 3445
rect 1150 3411 1184 3445
rect 1222 3411 1256 3445
rect 1078 3339 1112 3373
rect 1150 3339 1184 3373
rect 1222 3339 1256 3373
rect 1078 3267 1112 3301
rect 1150 3267 1184 3301
rect 1222 3267 1256 3301
rect 1078 3195 1112 3229
rect 1150 3195 1184 3229
rect 1222 3195 1256 3229
rect 1078 3123 1112 3157
rect 1150 3123 1184 3157
rect 1222 3123 1256 3157
rect 1078 3051 1112 3085
rect 1150 3051 1184 3085
rect 1222 3051 1256 3085
rect 1078 2979 1112 3013
rect 1150 2979 1184 3013
rect 1222 2979 1256 3013
rect 1078 2907 1112 2941
rect 1150 2907 1184 2941
rect 1222 2907 1256 2941
rect 1078 2835 1112 2869
rect 1150 2835 1184 2869
rect 1222 2835 1256 2869
rect 1078 2763 1112 2797
rect 1150 2763 1184 2797
rect 1222 2763 1256 2797
rect 1078 2691 1112 2725
rect 1150 2691 1184 2725
rect 1222 2691 1256 2725
rect 1078 2619 1112 2653
rect 1150 2619 1184 2653
rect 1222 2619 1256 2653
rect 1078 2547 1112 2581
rect 1150 2547 1184 2581
rect 1222 2547 1256 2581
rect 1078 2475 1112 2509
rect 1150 2475 1184 2509
rect 1222 2475 1256 2509
rect 1078 2403 1112 2437
rect 1150 2403 1184 2437
rect 1222 2403 1256 2437
rect 1078 2331 1112 2365
rect 1150 2331 1184 2365
rect 1222 2331 1256 2365
rect 1078 2259 1112 2293
rect 1150 2259 1184 2293
rect 1222 2259 1256 2293
rect 1078 2187 1112 2221
rect 1150 2187 1184 2221
rect 1222 2187 1256 2221
rect 1078 2115 1112 2149
rect 1150 2115 1184 2149
rect 1222 2115 1256 2149
rect 1078 2043 1112 2077
rect 1150 2043 1184 2077
rect 1222 2043 1256 2077
rect 1078 1971 1112 2005
rect 1150 1971 1184 2005
rect 1222 1971 1256 2005
rect 1078 1899 1112 1933
rect 1150 1899 1184 1933
rect 1222 1899 1256 1933
rect 1078 1827 1112 1861
rect 1150 1827 1184 1861
rect 1222 1827 1256 1861
rect 1078 1755 1112 1789
rect 1150 1755 1184 1789
rect 1222 1755 1256 1789
rect 1078 1683 1112 1717
rect 1150 1683 1184 1717
rect 1222 1683 1256 1717
rect 1078 1611 1112 1645
rect 1150 1611 1184 1645
rect 1222 1611 1256 1645
rect 1078 1539 1112 1573
rect 1150 1539 1184 1573
rect 1222 1539 1256 1573
rect 1078 1467 1112 1501
rect 1150 1467 1184 1501
rect 1222 1467 1256 1501
rect 1078 1395 1112 1429
rect 1150 1395 1184 1429
rect 1222 1395 1256 1429
rect 1078 1323 1112 1357
rect 1150 1323 1184 1357
rect 1222 1323 1256 1357
rect 1078 1251 1112 1285
rect 1150 1251 1184 1285
rect 1222 1251 1256 1285
rect 1078 1179 1112 1213
rect 1150 1179 1184 1213
rect 1222 1179 1256 1213
rect 1078 1107 1112 1141
rect 1150 1107 1184 1141
rect 1222 1107 1256 1141
rect 1078 1035 1112 1069
rect 1150 1035 1184 1069
rect 1222 1035 1256 1069
rect 1078 963 1112 997
rect 1150 963 1184 997
rect 1222 963 1256 997
rect 1078 891 1112 925
rect 1150 891 1184 925
rect 1222 891 1256 925
rect 1078 819 1112 853
rect 1150 819 1184 853
rect 1222 819 1256 853
rect 1078 747 1112 781
rect 1150 747 1184 781
rect 1222 747 1256 781
rect 1078 675 1112 709
rect 1150 675 1184 709
rect 1222 675 1256 709
rect 1078 603 1112 637
rect 1150 603 1184 637
rect 1222 603 1256 637
rect 1078 531 1112 565
rect 1150 531 1184 565
rect 1222 531 1256 565
rect 1078 459 1112 493
rect 1150 459 1184 493
rect 1222 459 1256 493
rect 1078 387 1112 421
rect 1150 387 1184 421
rect 1222 387 1256 421
rect 1078 315 1112 349
rect 1150 315 1184 349
rect 1222 315 1256 349
rect 1078 243 1112 277
rect 1150 243 1184 277
rect 1222 243 1256 277
rect 1078 171 1112 205
rect 1150 171 1184 205
rect 1222 171 1256 205
rect 1078 99 1112 133
rect 1150 99 1184 133
rect 1222 99 1256 133
<< nsubdiff >>
rect 1269 8053 1534 8076
rect 1269 8019 1313 8053
rect 1347 8019 1385 8053
rect 1419 8019 1457 8053
rect 1491 8019 1534 8053
rect 1269 7981 1534 8019
rect 1269 7947 1313 7981
rect 1347 7947 1385 7981
rect 1419 7947 1457 7981
rect 1491 7947 1534 7981
rect 1269 7909 1534 7947
rect 1269 7875 1313 7909
rect 1347 7875 1385 7909
rect 1419 7875 1457 7909
rect 1491 7875 1534 7909
rect 1269 7837 1534 7875
rect 1269 7803 1313 7837
rect 1347 7803 1385 7837
rect 1419 7803 1457 7837
rect 1491 7803 1534 7837
rect 1269 7765 1534 7803
rect 1269 7731 1313 7765
rect 1347 7731 1385 7765
rect 1419 7731 1457 7765
rect 1491 7731 1534 7765
rect 1269 7693 1534 7731
rect 1269 7659 1313 7693
rect 1347 7659 1385 7693
rect 1419 7659 1457 7693
rect 1491 7659 1534 7693
rect 1269 7621 1534 7659
rect 1269 7587 1313 7621
rect 1347 7587 1385 7621
rect 1419 7587 1457 7621
rect 1491 7587 1534 7621
rect 1269 7549 1534 7587
rect 1269 7515 1313 7549
rect 1347 7515 1385 7549
rect 1419 7515 1457 7549
rect 1491 7515 1534 7549
rect 1269 7477 1534 7515
rect 1269 7443 1313 7477
rect 1347 7443 1385 7477
rect 1419 7443 1457 7477
rect 1491 7443 1534 7477
rect 1269 7405 1534 7443
rect 1269 7371 1313 7405
rect 1347 7371 1385 7405
rect 1419 7371 1457 7405
rect 1491 7371 1534 7405
rect 1269 7333 1534 7371
rect 1269 7299 1313 7333
rect 1347 7299 1385 7333
rect 1419 7299 1457 7333
rect 1491 7299 1534 7333
rect 1269 7261 1534 7299
rect 1269 7227 1313 7261
rect 1347 7227 1385 7261
rect 1419 7227 1457 7261
rect 1491 7227 1534 7261
rect 1269 7189 1534 7227
rect 1269 7155 1313 7189
rect 1347 7155 1385 7189
rect 1419 7155 1457 7189
rect 1491 7155 1534 7189
rect 1269 7117 1534 7155
rect 1269 7083 1313 7117
rect 1347 7083 1385 7117
rect 1419 7083 1457 7117
rect 1491 7083 1534 7117
rect 1269 7045 1534 7083
rect 1269 7011 1313 7045
rect 1347 7011 1385 7045
rect 1419 7011 1457 7045
rect 1491 7011 1534 7045
rect 1269 6973 1534 7011
rect 1269 6939 1313 6973
rect 1347 6939 1385 6973
rect 1419 6939 1457 6973
rect 1491 6939 1534 6973
rect 1269 6901 1534 6939
rect 1269 6867 1313 6901
rect 1347 6867 1385 6901
rect 1419 6867 1457 6901
rect 1491 6867 1534 6901
rect 1269 6829 1534 6867
rect 1269 6795 1313 6829
rect 1347 6795 1385 6829
rect 1419 6795 1457 6829
rect 1491 6795 1534 6829
rect 1269 6757 1534 6795
rect 1269 6723 1313 6757
rect 1347 6723 1385 6757
rect 1419 6723 1457 6757
rect 1491 6723 1534 6757
rect 1269 6685 1534 6723
rect 1269 6651 1313 6685
rect 1347 6651 1385 6685
rect 1419 6651 1457 6685
rect 1491 6651 1534 6685
rect 1269 6613 1534 6651
rect 1269 6579 1313 6613
rect 1347 6579 1385 6613
rect 1419 6579 1457 6613
rect 1491 6579 1534 6613
rect 1269 6541 1534 6579
rect 1269 6507 1313 6541
rect 1347 6507 1385 6541
rect 1419 6507 1457 6541
rect 1491 6507 1534 6541
rect 1269 6469 1534 6507
rect 1269 6435 1313 6469
rect 1347 6435 1385 6469
rect 1419 6435 1457 6469
rect 1491 6435 1534 6469
rect 1269 6397 1534 6435
rect 1269 6363 1313 6397
rect 1347 6363 1385 6397
rect 1419 6363 1457 6397
rect 1491 6363 1534 6397
rect 1269 6325 1534 6363
rect 1269 6291 1313 6325
rect 1347 6291 1385 6325
rect 1419 6291 1457 6325
rect 1491 6291 1534 6325
rect 1269 6253 1534 6291
rect 1269 6219 1313 6253
rect 1347 6219 1385 6253
rect 1419 6219 1457 6253
rect 1491 6219 1534 6253
rect 1269 6181 1534 6219
rect 1269 6147 1313 6181
rect 1347 6147 1385 6181
rect 1419 6147 1457 6181
rect 1491 6147 1534 6181
rect 1269 6109 1534 6147
rect 1269 6075 1313 6109
rect 1347 6075 1385 6109
rect 1419 6075 1457 6109
rect 1491 6075 1534 6109
rect 1269 6037 1534 6075
rect 1269 6003 1313 6037
rect 1347 6003 1385 6037
rect 1419 6003 1457 6037
rect 1491 6003 1534 6037
rect 1269 5965 1534 6003
rect 1269 5931 1313 5965
rect 1347 5931 1385 5965
rect 1419 5931 1457 5965
rect 1491 5931 1534 5965
rect 1269 5893 1534 5931
rect 1269 5859 1313 5893
rect 1347 5859 1385 5893
rect 1419 5859 1457 5893
rect 1491 5859 1534 5893
rect 1269 5821 1534 5859
rect 1269 5787 1313 5821
rect 1347 5787 1385 5821
rect 1419 5787 1457 5821
rect 1491 5787 1534 5821
rect 1269 5749 1534 5787
rect 1269 5715 1313 5749
rect 1347 5715 1385 5749
rect 1419 5715 1457 5749
rect 1491 5715 1534 5749
rect 1269 5677 1534 5715
rect 1269 5643 1313 5677
rect 1347 5643 1385 5677
rect 1419 5643 1457 5677
rect 1491 5643 1534 5677
rect 1269 5605 1534 5643
rect 1269 5571 1313 5605
rect 1347 5571 1385 5605
rect 1419 5571 1457 5605
rect 1491 5571 1534 5605
rect 1269 5533 1534 5571
rect 1269 5499 1313 5533
rect 1347 5499 1385 5533
rect 1419 5499 1457 5533
rect 1491 5499 1534 5533
rect 1269 5461 1534 5499
rect 1269 5427 1313 5461
rect 1347 5427 1385 5461
rect 1419 5427 1457 5461
rect 1491 5427 1534 5461
rect 1269 5389 1534 5427
rect 1269 5355 1313 5389
rect 1347 5355 1385 5389
rect 1419 5355 1457 5389
rect 1491 5355 1534 5389
rect 1269 5317 1534 5355
rect 1269 5283 1313 5317
rect 1347 5283 1385 5317
rect 1419 5283 1457 5317
rect 1491 5283 1534 5317
rect 1269 5245 1534 5283
rect 1269 5211 1313 5245
rect 1347 5211 1385 5245
rect 1419 5211 1457 5245
rect 1491 5211 1534 5245
rect 1269 5173 1534 5211
rect 1269 5139 1313 5173
rect 1347 5139 1385 5173
rect 1419 5139 1457 5173
rect 1491 5139 1534 5173
rect 1269 5101 1534 5139
rect 1269 5067 1313 5101
rect 1347 5067 1385 5101
rect 1419 5067 1457 5101
rect 1491 5067 1534 5101
rect 1269 5029 1534 5067
rect 1269 4995 1313 5029
rect 1347 4995 1385 5029
rect 1419 4995 1457 5029
rect 1491 4995 1534 5029
rect 1269 4957 1534 4995
rect 1269 4923 1313 4957
rect 1347 4923 1385 4957
rect 1419 4923 1457 4957
rect 1491 4923 1534 4957
rect 1269 4885 1534 4923
rect 1269 4851 1313 4885
rect 1347 4851 1385 4885
rect 1419 4851 1457 4885
rect 1491 4851 1534 4885
rect 1269 4813 1534 4851
rect 1269 4779 1313 4813
rect 1347 4779 1385 4813
rect 1419 4779 1457 4813
rect 1491 4779 1534 4813
rect 1269 4741 1534 4779
rect 1269 4707 1313 4741
rect 1347 4707 1385 4741
rect 1419 4707 1457 4741
rect 1491 4707 1534 4741
rect 1269 4669 1534 4707
rect 1269 4635 1313 4669
rect 1347 4635 1385 4669
rect 1419 4635 1457 4669
rect 1491 4635 1534 4669
rect 1269 4597 1534 4635
rect 1269 4563 1313 4597
rect 1347 4563 1385 4597
rect 1419 4563 1457 4597
rect 1491 4563 1534 4597
rect 1269 4525 1534 4563
rect 1269 4491 1313 4525
rect 1347 4491 1385 4525
rect 1419 4491 1457 4525
rect 1491 4491 1534 4525
rect 1269 4453 1534 4491
rect 1269 4419 1313 4453
rect 1347 4419 1385 4453
rect 1419 4419 1457 4453
rect 1491 4419 1534 4453
rect 1269 4381 1534 4419
rect 1269 4347 1313 4381
rect 1347 4347 1385 4381
rect 1419 4347 1457 4381
rect 1491 4347 1534 4381
rect 1269 4309 1534 4347
rect 1269 4275 1313 4309
rect 1347 4275 1385 4309
rect 1419 4275 1457 4309
rect 1491 4275 1534 4309
rect 1269 4237 1534 4275
rect 1269 4203 1313 4237
rect 1347 4203 1385 4237
rect 1419 4203 1457 4237
rect 1491 4203 1534 4237
rect 1269 4165 1534 4203
rect 1269 4131 1313 4165
rect 1347 4131 1385 4165
rect 1419 4131 1457 4165
rect 1491 4131 1534 4165
rect 1269 4093 1534 4131
rect 1269 4059 1313 4093
rect 1347 4059 1385 4093
rect 1419 4059 1457 4093
rect 1491 4059 1534 4093
rect 1269 4021 1534 4059
rect 1269 3987 1313 4021
rect 1347 3987 1385 4021
rect 1419 3987 1457 4021
rect 1491 3987 1534 4021
rect 1269 3949 1534 3987
rect 1269 3915 1313 3949
rect 1347 3915 1385 3949
rect 1419 3915 1457 3949
rect 1491 3915 1534 3949
rect 1269 3877 1534 3915
rect 1269 3843 1313 3877
rect 1347 3843 1385 3877
rect 1419 3843 1457 3877
rect 1491 3843 1534 3877
rect 1269 3805 1534 3843
rect 1269 3771 1313 3805
rect 1347 3771 1385 3805
rect 1419 3771 1457 3805
rect 1491 3771 1534 3805
rect 1269 3733 1534 3771
rect 1269 3699 1313 3733
rect 1347 3699 1385 3733
rect 1419 3699 1457 3733
rect 1491 3699 1534 3733
rect 1269 3661 1534 3699
rect 1269 3627 1313 3661
rect 1347 3627 1385 3661
rect 1419 3627 1457 3661
rect 1491 3627 1534 3661
rect 1269 3589 1534 3627
rect 1269 3555 1313 3589
rect 1347 3555 1385 3589
rect 1419 3555 1457 3589
rect 1491 3555 1534 3589
rect 1269 3517 1534 3555
rect 1269 3483 1313 3517
rect 1347 3483 1385 3517
rect 1419 3483 1457 3517
rect 1491 3483 1534 3517
rect 1269 3445 1534 3483
rect 1269 3411 1313 3445
rect 1347 3411 1385 3445
rect 1419 3411 1457 3445
rect 1491 3411 1534 3445
rect 1269 3373 1534 3411
rect 1269 3339 1313 3373
rect 1347 3339 1385 3373
rect 1419 3339 1457 3373
rect 1491 3339 1534 3373
rect 1269 3301 1534 3339
rect 1269 3267 1313 3301
rect 1347 3267 1385 3301
rect 1419 3267 1457 3301
rect 1491 3267 1534 3301
rect 1269 3229 1534 3267
rect 1269 3195 1313 3229
rect 1347 3195 1385 3229
rect 1419 3195 1457 3229
rect 1491 3195 1534 3229
rect 1269 3157 1534 3195
rect 1269 3123 1313 3157
rect 1347 3123 1385 3157
rect 1419 3123 1457 3157
rect 1491 3123 1534 3157
rect 1269 3085 1534 3123
rect 1269 3051 1313 3085
rect 1347 3051 1385 3085
rect 1419 3051 1457 3085
rect 1491 3051 1534 3085
rect 1269 3013 1534 3051
rect 1269 2979 1313 3013
rect 1347 2979 1385 3013
rect 1419 2979 1457 3013
rect 1491 2979 1534 3013
rect 1269 2941 1534 2979
rect 1269 2907 1313 2941
rect 1347 2907 1385 2941
rect 1419 2907 1457 2941
rect 1491 2907 1534 2941
rect 1269 2869 1534 2907
rect 1269 2835 1313 2869
rect 1347 2835 1385 2869
rect 1419 2835 1457 2869
rect 1491 2835 1534 2869
rect 1269 2797 1534 2835
rect 1269 2763 1313 2797
rect 1347 2763 1385 2797
rect 1419 2763 1457 2797
rect 1491 2763 1534 2797
rect 1269 2725 1534 2763
rect 1269 2691 1313 2725
rect 1347 2691 1385 2725
rect 1419 2691 1457 2725
rect 1491 2691 1534 2725
rect 1269 2653 1534 2691
rect 1269 2619 1313 2653
rect 1347 2619 1385 2653
rect 1419 2619 1457 2653
rect 1491 2619 1534 2653
rect 1269 2581 1534 2619
rect 1269 2547 1313 2581
rect 1347 2547 1385 2581
rect 1419 2547 1457 2581
rect 1491 2547 1534 2581
rect 1269 2509 1534 2547
rect 1269 2475 1313 2509
rect 1347 2475 1385 2509
rect 1419 2475 1457 2509
rect 1491 2475 1534 2509
rect 1269 2437 1534 2475
rect 1269 2403 1313 2437
rect 1347 2403 1385 2437
rect 1419 2403 1457 2437
rect 1491 2403 1534 2437
rect 1269 2365 1534 2403
rect 1269 2331 1313 2365
rect 1347 2331 1385 2365
rect 1419 2331 1457 2365
rect 1491 2331 1534 2365
rect 1269 2293 1534 2331
rect 1269 2259 1313 2293
rect 1347 2259 1385 2293
rect 1419 2259 1457 2293
rect 1491 2259 1534 2293
rect 1269 2221 1534 2259
rect 1269 2187 1313 2221
rect 1347 2187 1385 2221
rect 1419 2187 1457 2221
rect 1491 2187 1534 2221
rect 1269 2149 1534 2187
rect 1269 2115 1313 2149
rect 1347 2115 1385 2149
rect 1419 2115 1457 2149
rect 1491 2115 1534 2149
rect 1269 2077 1534 2115
rect 1269 2043 1313 2077
rect 1347 2043 1385 2077
rect 1419 2043 1457 2077
rect 1491 2043 1534 2077
rect 1269 2005 1534 2043
rect 1269 1971 1313 2005
rect 1347 1971 1385 2005
rect 1419 1971 1457 2005
rect 1491 1971 1534 2005
rect 1269 1933 1534 1971
rect 1269 1899 1313 1933
rect 1347 1899 1385 1933
rect 1419 1899 1457 1933
rect 1491 1899 1534 1933
rect 1269 1861 1534 1899
rect 1269 1827 1313 1861
rect 1347 1827 1385 1861
rect 1419 1827 1457 1861
rect 1491 1827 1534 1861
rect 1269 1789 1534 1827
rect 1269 1755 1313 1789
rect 1347 1755 1385 1789
rect 1419 1755 1457 1789
rect 1491 1755 1534 1789
rect 1269 1717 1534 1755
rect 1269 1683 1313 1717
rect 1347 1683 1385 1717
rect 1419 1683 1457 1717
rect 1491 1683 1534 1717
rect 1269 1645 1534 1683
rect 1269 1611 1313 1645
rect 1347 1611 1385 1645
rect 1419 1611 1457 1645
rect 1491 1611 1534 1645
rect 1269 1573 1534 1611
rect 1269 1539 1313 1573
rect 1347 1539 1385 1573
rect 1419 1539 1457 1573
rect 1491 1539 1534 1573
rect 1269 1501 1534 1539
rect 1269 1467 1313 1501
rect 1347 1467 1385 1501
rect 1419 1467 1457 1501
rect 1491 1467 1534 1501
rect 1269 1429 1534 1467
rect 1269 1395 1313 1429
rect 1347 1395 1385 1429
rect 1419 1395 1457 1429
rect 1491 1395 1534 1429
rect 1269 1357 1534 1395
rect 1269 1323 1313 1357
rect 1347 1323 1385 1357
rect 1419 1323 1457 1357
rect 1491 1323 1534 1357
rect 1269 1285 1534 1323
rect 1269 1251 1313 1285
rect 1347 1251 1385 1285
rect 1419 1251 1457 1285
rect 1491 1251 1534 1285
rect 1269 1213 1534 1251
rect 1269 1179 1313 1213
rect 1347 1179 1385 1213
rect 1419 1179 1457 1213
rect 1491 1179 1534 1213
rect 1269 1141 1534 1179
rect 1269 1107 1313 1141
rect 1347 1107 1385 1141
rect 1419 1107 1457 1141
rect 1491 1107 1534 1141
rect 1269 1069 1534 1107
rect 1269 1035 1313 1069
rect 1347 1035 1385 1069
rect 1419 1035 1457 1069
rect 1491 1035 1534 1069
rect 1269 997 1534 1035
rect 1269 963 1313 997
rect 1347 963 1385 997
rect 1419 963 1457 997
rect 1491 963 1534 997
rect 1269 925 1534 963
rect 1269 891 1313 925
rect 1347 891 1385 925
rect 1419 891 1457 925
rect 1491 891 1534 925
rect 1269 853 1534 891
rect 1269 819 1313 853
rect 1347 819 1385 853
rect 1419 819 1457 853
rect 1491 819 1534 853
rect 1269 781 1534 819
rect 1269 747 1313 781
rect 1347 747 1385 781
rect 1419 747 1457 781
rect 1491 747 1534 781
rect 1269 709 1534 747
rect 1269 675 1313 709
rect 1347 675 1385 709
rect 1419 675 1457 709
rect 1491 675 1534 709
rect 1269 637 1534 675
rect 1269 603 1313 637
rect 1347 603 1385 637
rect 1419 603 1457 637
rect 1491 603 1534 637
rect 1269 565 1534 603
rect 1269 531 1313 565
rect 1347 531 1385 565
rect 1419 531 1457 565
rect 1491 531 1534 565
rect 1269 493 1534 531
rect 1269 459 1313 493
rect 1347 459 1385 493
rect 1419 459 1457 493
rect 1491 459 1534 493
rect 1269 421 1534 459
rect 1269 387 1313 421
rect 1347 387 1385 421
rect 1419 387 1457 421
rect 1491 387 1534 421
rect 1269 349 1534 387
rect 1269 315 1313 349
rect 1347 315 1385 349
rect 1419 315 1457 349
rect 1491 315 1534 349
rect 1269 277 1534 315
rect 1269 243 1313 277
rect 1347 243 1385 277
rect 1419 243 1457 277
rect 1491 243 1534 277
rect 1269 205 1534 243
rect 1269 171 1313 205
rect 1347 171 1385 205
rect 1419 171 1457 205
rect 1491 171 1534 205
rect 1269 133 1534 171
rect 1269 99 1313 133
rect 1347 99 1385 133
rect 1419 99 1457 133
rect 1491 99 1534 133
rect 1269 76 1534 99
<< nsubdiffcont >>
rect 1313 8019 1347 8053
rect 1385 8019 1419 8053
rect 1457 8019 1491 8053
rect 1313 7947 1347 7981
rect 1385 7947 1419 7981
rect 1457 7947 1491 7981
rect 1313 7875 1347 7909
rect 1385 7875 1419 7909
rect 1457 7875 1491 7909
rect 1313 7803 1347 7837
rect 1385 7803 1419 7837
rect 1457 7803 1491 7837
rect 1313 7731 1347 7765
rect 1385 7731 1419 7765
rect 1457 7731 1491 7765
rect 1313 7659 1347 7693
rect 1385 7659 1419 7693
rect 1457 7659 1491 7693
rect 1313 7587 1347 7621
rect 1385 7587 1419 7621
rect 1457 7587 1491 7621
rect 1313 7515 1347 7549
rect 1385 7515 1419 7549
rect 1457 7515 1491 7549
rect 1313 7443 1347 7477
rect 1385 7443 1419 7477
rect 1457 7443 1491 7477
rect 1313 7371 1347 7405
rect 1385 7371 1419 7405
rect 1457 7371 1491 7405
rect 1313 7299 1347 7333
rect 1385 7299 1419 7333
rect 1457 7299 1491 7333
rect 1313 7227 1347 7261
rect 1385 7227 1419 7261
rect 1457 7227 1491 7261
rect 1313 7155 1347 7189
rect 1385 7155 1419 7189
rect 1457 7155 1491 7189
rect 1313 7083 1347 7117
rect 1385 7083 1419 7117
rect 1457 7083 1491 7117
rect 1313 7011 1347 7045
rect 1385 7011 1419 7045
rect 1457 7011 1491 7045
rect 1313 6939 1347 6973
rect 1385 6939 1419 6973
rect 1457 6939 1491 6973
rect 1313 6867 1347 6901
rect 1385 6867 1419 6901
rect 1457 6867 1491 6901
rect 1313 6795 1347 6829
rect 1385 6795 1419 6829
rect 1457 6795 1491 6829
rect 1313 6723 1347 6757
rect 1385 6723 1419 6757
rect 1457 6723 1491 6757
rect 1313 6651 1347 6685
rect 1385 6651 1419 6685
rect 1457 6651 1491 6685
rect 1313 6579 1347 6613
rect 1385 6579 1419 6613
rect 1457 6579 1491 6613
rect 1313 6507 1347 6541
rect 1385 6507 1419 6541
rect 1457 6507 1491 6541
rect 1313 6435 1347 6469
rect 1385 6435 1419 6469
rect 1457 6435 1491 6469
rect 1313 6363 1347 6397
rect 1385 6363 1419 6397
rect 1457 6363 1491 6397
rect 1313 6291 1347 6325
rect 1385 6291 1419 6325
rect 1457 6291 1491 6325
rect 1313 6219 1347 6253
rect 1385 6219 1419 6253
rect 1457 6219 1491 6253
rect 1313 6147 1347 6181
rect 1385 6147 1419 6181
rect 1457 6147 1491 6181
rect 1313 6075 1347 6109
rect 1385 6075 1419 6109
rect 1457 6075 1491 6109
rect 1313 6003 1347 6037
rect 1385 6003 1419 6037
rect 1457 6003 1491 6037
rect 1313 5931 1347 5965
rect 1385 5931 1419 5965
rect 1457 5931 1491 5965
rect 1313 5859 1347 5893
rect 1385 5859 1419 5893
rect 1457 5859 1491 5893
rect 1313 5787 1347 5821
rect 1385 5787 1419 5821
rect 1457 5787 1491 5821
rect 1313 5715 1347 5749
rect 1385 5715 1419 5749
rect 1457 5715 1491 5749
rect 1313 5643 1347 5677
rect 1385 5643 1419 5677
rect 1457 5643 1491 5677
rect 1313 5571 1347 5605
rect 1385 5571 1419 5605
rect 1457 5571 1491 5605
rect 1313 5499 1347 5533
rect 1385 5499 1419 5533
rect 1457 5499 1491 5533
rect 1313 5427 1347 5461
rect 1385 5427 1419 5461
rect 1457 5427 1491 5461
rect 1313 5355 1347 5389
rect 1385 5355 1419 5389
rect 1457 5355 1491 5389
rect 1313 5283 1347 5317
rect 1385 5283 1419 5317
rect 1457 5283 1491 5317
rect 1313 5211 1347 5245
rect 1385 5211 1419 5245
rect 1457 5211 1491 5245
rect 1313 5139 1347 5173
rect 1385 5139 1419 5173
rect 1457 5139 1491 5173
rect 1313 5067 1347 5101
rect 1385 5067 1419 5101
rect 1457 5067 1491 5101
rect 1313 4995 1347 5029
rect 1385 4995 1419 5029
rect 1457 4995 1491 5029
rect 1313 4923 1347 4957
rect 1385 4923 1419 4957
rect 1457 4923 1491 4957
rect 1313 4851 1347 4885
rect 1385 4851 1419 4885
rect 1457 4851 1491 4885
rect 1313 4779 1347 4813
rect 1385 4779 1419 4813
rect 1457 4779 1491 4813
rect 1313 4707 1347 4741
rect 1385 4707 1419 4741
rect 1457 4707 1491 4741
rect 1313 4635 1347 4669
rect 1385 4635 1419 4669
rect 1457 4635 1491 4669
rect 1313 4563 1347 4597
rect 1385 4563 1419 4597
rect 1457 4563 1491 4597
rect 1313 4491 1347 4525
rect 1385 4491 1419 4525
rect 1457 4491 1491 4525
rect 1313 4419 1347 4453
rect 1385 4419 1419 4453
rect 1457 4419 1491 4453
rect 1313 4347 1347 4381
rect 1385 4347 1419 4381
rect 1457 4347 1491 4381
rect 1313 4275 1347 4309
rect 1385 4275 1419 4309
rect 1457 4275 1491 4309
rect 1313 4203 1347 4237
rect 1385 4203 1419 4237
rect 1457 4203 1491 4237
rect 1313 4131 1347 4165
rect 1385 4131 1419 4165
rect 1457 4131 1491 4165
rect 1313 4059 1347 4093
rect 1385 4059 1419 4093
rect 1457 4059 1491 4093
rect 1313 3987 1347 4021
rect 1385 3987 1419 4021
rect 1457 3987 1491 4021
rect 1313 3915 1347 3949
rect 1385 3915 1419 3949
rect 1457 3915 1491 3949
rect 1313 3843 1347 3877
rect 1385 3843 1419 3877
rect 1457 3843 1491 3877
rect 1313 3771 1347 3805
rect 1385 3771 1419 3805
rect 1457 3771 1491 3805
rect 1313 3699 1347 3733
rect 1385 3699 1419 3733
rect 1457 3699 1491 3733
rect 1313 3627 1347 3661
rect 1385 3627 1419 3661
rect 1457 3627 1491 3661
rect 1313 3555 1347 3589
rect 1385 3555 1419 3589
rect 1457 3555 1491 3589
rect 1313 3483 1347 3517
rect 1385 3483 1419 3517
rect 1457 3483 1491 3517
rect 1313 3411 1347 3445
rect 1385 3411 1419 3445
rect 1457 3411 1491 3445
rect 1313 3339 1347 3373
rect 1385 3339 1419 3373
rect 1457 3339 1491 3373
rect 1313 3267 1347 3301
rect 1385 3267 1419 3301
rect 1457 3267 1491 3301
rect 1313 3195 1347 3229
rect 1385 3195 1419 3229
rect 1457 3195 1491 3229
rect 1313 3123 1347 3157
rect 1385 3123 1419 3157
rect 1457 3123 1491 3157
rect 1313 3051 1347 3085
rect 1385 3051 1419 3085
rect 1457 3051 1491 3085
rect 1313 2979 1347 3013
rect 1385 2979 1419 3013
rect 1457 2979 1491 3013
rect 1313 2907 1347 2941
rect 1385 2907 1419 2941
rect 1457 2907 1491 2941
rect 1313 2835 1347 2869
rect 1385 2835 1419 2869
rect 1457 2835 1491 2869
rect 1313 2763 1347 2797
rect 1385 2763 1419 2797
rect 1457 2763 1491 2797
rect 1313 2691 1347 2725
rect 1385 2691 1419 2725
rect 1457 2691 1491 2725
rect 1313 2619 1347 2653
rect 1385 2619 1419 2653
rect 1457 2619 1491 2653
rect 1313 2547 1347 2581
rect 1385 2547 1419 2581
rect 1457 2547 1491 2581
rect 1313 2475 1347 2509
rect 1385 2475 1419 2509
rect 1457 2475 1491 2509
rect 1313 2403 1347 2437
rect 1385 2403 1419 2437
rect 1457 2403 1491 2437
rect 1313 2331 1347 2365
rect 1385 2331 1419 2365
rect 1457 2331 1491 2365
rect 1313 2259 1347 2293
rect 1385 2259 1419 2293
rect 1457 2259 1491 2293
rect 1313 2187 1347 2221
rect 1385 2187 1419 2221
rect 1457 2187 1491 2221
rect 1313 2115 1347 2149
rect 1385 2115 1419 2149
rect 1457 2115 1491 2149
rect 1313 2043 1347 2077
rect 1385 2043 1419 2077
rect 1457 2043 1491 2077
rect 1313 1971 1347 2005
rect 1385 1971 1419 2005
rect 1457 1971 1491 2005
rect 1313 1899 1347 1933
rect 1385 1899 1419 1933
rect 1457 1899 1491 1933
rect 1313 1827 1347 1861
rect 1385 1827 1419 1861
rect 1457 1827 1491 1861
rect 1313 1755 1347 1789
rect 1385 1755 1419 1789
rect 1457 1755 1491 1789
rect 1313 1683 1347 1717
rect 1385 1683 1419 1717
rect 1457 1683 1491 1717
rect 1313 1611 1347 1645
rect 1385 1611 1419 1645
rect 1457 1611 1491 1645
rect 1313 1539 1347 1573
rect 1385 1539 1419 1573
rect 1457 1539 1491 1573
rect 1313 1467 1347 1501
rect 1385 1467 1419 1501
rect 1457 1467 1491 1501
rect 1313 1395 1347 1429
rect 1385 1395 1419 1429
rect 1457 1395 1491 1429
rect 1313 1323 1347 1357
rect 1385 1323 1419 1357
rect 1457 1323 1491 1357
rect 1313 1251 1347 1285
rect 1385 1251 1419 1285
rect 1457 1251 1491 1285
rect 1313 1179 1347 1213
rect 1385 1179 1419 1213
rect 1457 1179 1491 1213
rect 1313 1107 1347 1141
rect 1385 1107 1419 1141
rect 1457 1107 1491 1141
rect 1313 1035 1347 1069
rect 1385 1035 1419 1069
rect 1457 1035 1491 1069
rect 1313 963 1347 997
rect 1385 963 1419 997
rect 1457 963 1491 997
rect 1313 891 1347 925
rect 1385 891 1419 925
rect 1457 891 1491 925
rect 1313 819 1347 853
rect 1385 819 1419 853
rect 1457 819 1491 853
rect 1313 747 1347 781
rect 1385 747 1419 781
rect 1457 747 1491 781
rect 1313 675 1347 709
rect 1385 675 1419 709
rect 1457 675 1491 709
rect 1313 603 1347 637
rect 1385 603 1419 637
rect 1457 603 1491 637
rect 1313 531 1347 565
rect 1385 531 1419 565
rect 1457 531 1491 565
rect 1313 459 1347 493
rect 1385 459 1419 493
rect 1457 459 1491 493
rect 1313 387 1347 421
rect 1385 387 1419 421
rect 1457 387 1491 421
rect 1313 315 1347 349
rect 1385 315 1419 349
rect 1457 315 1491 349
rect 1313 243 1347 277
rect 1385 243 1419 277
rect 1457 243 1491 277
rect 1313 171 1347 205
rect 1385 171 1419 205
rect 1457 171 1491 205
rect 1313 99 1347 133
rect 1385 99 1419 133
rect 1457 99 1491 133
<< poly >>
rect 265 8166 1065 8182
rect 265 8132 288 8166
rect 322 8132 360 8166
rect 394 8132 432 8166
rect 466 8132 504 8166
rect 538 8132 576 8166
rect 610 8132 648 8166
rect 682 8132 720 8166
rect 754 8132 792 8166
rect 826 8132 864 8166
rect 898 8132 936 8166
rect 970 8132 1008 8166
rect 1042 8132 1065 8166
rect 265 8076 1065 8132
rect 265 36 1065 76
<< polycont >>
rect 288 8132 322 8166
rect 360 8132 394 8166
rect 432 8132 466 8166
rect 504 8132 538 8166
rect 576 8132 610 8166
rect 648 8132 682 8166
rect 720 8132 754 8166
rect 792 8132 826 8166
rect 864 8132 898 8166
rect 936 8132 970 8166
rect 1008 8132 1042 8166
<< locali >>
rect 272 8132 288 8166
rect 322 8132 360 8166
rect 394 8132 432 8166
rect 466 8132 504 8166
rect 538 8132 576 8166
rect 610 8132 648 8166
rect 682 8132 720 8166
rect 754 8132 792 8166
rect 826 8132 864 8166
rect 898 8132 936 8166
rect 970 8132 1008 8166
rect 1042 8132 1058 8166
rect 74 8053 252 8069
rect 74 83 252 99
rect 1078 8053 1256 8069
rect 1078 83 1256 99
rect 1313 8053 1491 8069
rect 1347 8019 1385 8053
rect 1419 8019 1457 8053
rect 1313 7981 1491 8019
rect 1347 7947 1385 7981
rect 1419 7947 1457 7981
rect 1313 7909 1491 7947
rect 1347 7875 1385 7909
rect 1419 7875 1457 7909
rect 1313 7837 1491 7875
rect 1347 7803 1385 7837
rect 1419 7803 1457 7837
rect 1313 7765 1491 7803
rect 1347 7731 1385 7765
rect 1419 7731 1457 7765
rect 1313 7693 1491 7731
rect 1347 7659 1385 7693
rect 1419 7659 1457 7693
rect 1313 7621 1491 7659
rect 1347 7587 1385 7621
rect 1419 7587 1457 7621
rect 1313 7549 1491 7587
rect 1347 7515 1385 7549
rect 1419 7515 1457 7549
rect 1313 7477 1491 7515
rect 1347 7443 1385 7477
rect 1419 7443 1457 7477
rect 1313 7405 1491 7443
rect 1347 7371 1385 7405
rect 1419 7371 1457 7405
rect 1313 7333 1491 7371
rect 1347 7299 1385 7333
rect 1419 7299 1457 7333
rect 1313 7261 1491 7299
rect 1347 7227 1385 7261
rect 1419 7227 1457 7261
rect 1313 7189 1491 7227
rect 1347 7155 1385 7189
rect 1419 7155 1457 7189
rect 1313 7117 1491 7155
rect 1347 7083 1385 7117
rect 1419 7083 1457 7117
rect 1313 7045 1491 7083
rect 1347 7011 1385 7045
rect 1419 7011 1457 7045
rect 1313 6973 1491 7011
rect 1347 6939 1385 6973
rect 1419 6939 1457 6973
rect 1313 6901 1491 6939
rect 1347 6867 1385 6901
rect 1419 6867 1457 6901
rect 1313 6829 1491 6867
rect 1347 6795 1385 6829
rect 1419 6795 1457 6829
rect 1313 6757 1491 6795
rect 1347 6723 1385 6757
rect 1419 6723 1457 6757
rect 1313 6685 1491 6723
rect 1347 6651 1385 6685
rect 1419 6651 1457 6685
rect 1313 6613 1491 6651
rect 1347 6579 1385 6613
rect 1419 6579 1457 6613
rect 1313 6541 1491 6579
rect 1347 6507 1385 6541
rect 1419 6507 1457 6541
rect 1313 6469 1491 6507
rect 1347 6435 1385 6469
rect 1419 6435 1457 6469
rect 1313 6397 1491 6435
rect 1347 6363 1385 6397
rect 1419 6363 1457 6397
rect 1313 6325 1491 6363
rect 1347 6291 1385 6325
rect 1419 6291 1457 6325
rect 1313 6253 1491 6291
rect 1347 6219 1385 6253
rect 1419 6219 1457 6253
rect 1313 6181 1491 6219
rect 1347 6147 1385 6181
rect 1419 6147 1457 6181
rect 1313 6109 1491 6147
rect 1347 6075 1385 6109
rect 1419 6075 1457 6109
rect 1313 6037 1491 6075
rect 1347 6003 1385 6037
rect 1419 6003 1457 6037
rect 1313 5965 1491 6003
rect 1347 5931 1385 5965
rect 1419 5931 1457 5965
rect 1313 5893 1491 5931
rect 1347 5859 1385 5893
rect 1419 5859 1457 5893
rect 1313 5821 1491 5859
rect 1347 5787 1385 5821
rect 1419 5787 1457 5821
rect 1313 5749 1491 5787
rect 1347 5715 1385 5749
rect 1419 5715 1457 5749
rect 1313 5677 1491 5715
rect 1347 5643 1385 5677
rect 1419 5643 1457 5677
rect 1313 5605 1491 5643
rect 1347 5571 1385 5605
rect 1419 5571 1457 5605
rect 1313 5533 1491 5571
rect 1347 5499 1385 5533
rect 1419 5499 1457 5533
rect 1313 5461 1491 5499
rect 1347 5427 1385 5461
rect 1419 5427 1457 5461
rect 1313 5389 1491 5427
rect 1347 5355 1385 5389
rect 1419 5355 1457 5389
rect 1313 5317 1491 5355
rect 1347 5283 1385 5317
rect 1419 5283 1457 5317
rect 1313 5245 1491 5283
rect 1347 5211 1385 5245
rect 1419 5211 1457 5245
rect 1313 5173 1491 5211
rect 1347 5139 1385 5173
rect 1419 5139 1457 5173
rect 1313 5101 1491 5139
rect 1347 5067 1385 5101
rect 1419 5067 1457 5101
rect 1313 5029 1491 5067
rect 1347 4995 1385 5029
rect 1419 4995 1457 5029
rect 1313 4957 1491 4995
rect 1347 4923 1385 4957
rect 1419 4923 1457 4957
rect 1313 4885 1491 4923
rect 1347 4851 1385 4885
rect 1419 4851 1457 4885
rect 1313 4813 1491 4851
rect 1347 4779 1385 4813
rect 1419 4779 1457 4813
rect 1313 4741 1491 4779
rect 1347 4707 1385 4741
rect 1419 4707 1457 4741
rect 1313 4669 1491 4707
rect 1347 4635 1385 4669
rect 1419 4635 1457 4669
rect 1313 4597 1491 4635
rect 1347 4563 1385 4597
rect 1419 4563 1457 4597
rect 1313 4525 1491 4563
rect 1347 4491 1385 4525
rect 1419 4491 1457 4525
rect 1313 4453 1491 4491
rect 1347 4419 1385 4453
rect 1419 4419 1457 4453
rect 1313 4381 1491 4419
rect 1347 4347 1385 4381
rect 1419 4347 1457 4381
rect 1313 4309 1491 4347
rect 1347 4275 1385 4309
rect 1419 4275 1457 4309
rect 1313 4237 1491 4275
rect 1347 4203 1385 4237
rect 1419 4203 1457 4237
rect 1313 4165 1491 4203
rect 1347 4131 1385 4165
rect 1419 4131 1457 4165
rect 1313 4093 1491 4131
rect 1347 4059 1385 4093
rect 1419 4059 1457 4093
rect 1313 4021 1491 4059
rect 1347 3987 1385 4021
rect 1419 3987 1457 4021
rect 1313 3949 1491 3987
rect 1347 3915 1385 3949
rect 1419 3915 1457 3949
rect 1313 3877 1491 3915
rect 1347 3843 1385 3877
rect 1419 3843 1457 3877
rect 1313 3805 1491 3843
rect 1347 3771 1385 3805
rect 1419 3771 1457 3805
rect 1313 3733 1491 3771
rect 1347 3699 1385 3733
rect 1419 3699 1457 3733
rect 1313 3661 1491 3699
rect 1347 3627 1385 3661
rect 1419 3627 1457 3661
rect 1313 3589 1491 3627
rect 1347 3555 1385 3589
rect 1419 3555 1457 3589
rect 1313 3517 1491 3555
rect 1347 3483 1385 3517
rect 1419 3483 1457 3517
rect 1313 3445 1491 3483
rect 1347 3411 1385 3445
rect 1419 3411 1457 3445
rect 1313 3373 1491 3411
rect 1347 3339 1385 3373
rect 1419 3339 1457 3373
rect 1313 3301 1491 3339
rect 1347 3267 1385 3301
rect 1419 3267 1457 3301
rect 1313 3229 1491 3267
rect 1347 3195 1385 3229
rect 1419 3195 1457 3229
rect 1313 3157 1491 3195
rect 1347 3123 1385 3157
rect 1419 3123 1457 3157
rect 1313 3085 1491 3123
rect 1347 3051 1385 3085
rect 1419 3051 1457 3085
rect 1313 3013 1491 3051
rect 1347 2979 1385 3013
rect 1419 2979 1457 3013
rect 1313 2941 1491 2979
rect 1347 2907 1385 2941
rect 1419 2907 1457 2941
rect 1313 2869 1491 2907
rect 1347 2835 1385 2869
rect 1419 2835 1457 2869
rect 1313 2797 1491 2835
rect 1347 2763 1385 2797
rect 1419 2763 1457 2797
rect 1313 2725 1491 2763
rect 1347 2691 1385 2725
rect 1419 2691 1457 2725
rect 1313 2653 1491 2691
rect 1347 2619 1385 2653
rect 1419 2619 1457 2653
rect 1313 2581 1491 2619
rect 1347 2547 1385 2581
rect 1419 2547 1457 2581
rect 1313 2509 1491 2547
rect 1347 2475 1385 2509
rect 1419 2475 1457 2509
rect 1313 2437 1491 2475
rect 1347 2403 1385 2437
rect 1419 2403 1457 2437
rect 1313 2365 1491 2403
rect 1347 2331 1385 2365
rect 1419 2331 1457 2365
rect 1313 2293 1491 2331
rect 1347 2259 1385 2293
rect 1419 2259 1457 2293
rect 1313 2221 1491 2259
rect 1347 2187 1385 2221
rect 1419 2187 1457 2221
rect 1313 2149 1491 2187
rect 1347 2115 1385 2149
rect 1419 2115 1457 2149
rect 1313 2077 1491 2115
rect 1347 2043 1385 2077
rect 1419 2043 1457 2077
rect 1313 2005 1491 2043
rect 1347 1971 1385 2005
rect 1419 1971 1457 2005
rect 1313 1933 1491 1971
rect 1347 1899 1385 1933
rect 1419 1899 1457 1933
rect 1313 1861 1491 1899
rect 1347 1827 1385 1861
rect 1419 1827 1457 1861
rect 1313 1789 1491 1827
rect 1347 1755 1385 1789
rect 1419 1755 1457 1789
rect 1313 1717 1491 1755
rect 1347 1683 1385 1717
rect 1419 1683 1457 1717
rect 1313 1645 1491 1683
rect 1347 1611 1385 1645
rect 1419 1611 1457 1645
rect 1313 1573 1491 1611
rect 1347 1539 1385 1573
rect 1419 1539 1457 1573
rect 1313 1501 1491 1539
rect 1347 1467 1385 1501
rect 1419 1467 1457 1501
rect 1313 1429 1491 1467
rect 1347 1395 1385 1429
rect 1419 1395 1457 1429
rect 1313 1357 1491 1395
rect 1347 1323 1385 1357
rect 1419 1323 1457 1357
rect 1313 1285 1491 1323
rect 1347 1251 1385 1285
rect 1419 1251 1457 1285
rect 1313 1213 1491 1251
rect 1347 1179 1385 1213
rect 1419 1179 1457 1213
rect 1313 1141 1491 1179
rect 1347 1107 1385 1141
rect 1419 1107 1457 1141
rect 1313 1069 1491 1107
rect 1347 1035 1385 1069
rect 1419 1035 1457 1069
rect 1313 997 1491 1035
rect 1347 963 1385 997
rect 1419 963 1457 997
rect 1313 925 1491 963
rect 1347 891 1385 925
rect 1419 891 1457 925
rect 1313 853 1491 891
rect 1347 819 1385 853
rect 1419 819 1457 853
rect 1313 781 1491 819
rect 1347 747 1385 781
rect 1419 747 1457 781
rect 1313 709 1491 747
rect 1347 675 1385 709
rect 1419 675 1457 709
rect 1313 637 1491 675
rect 1347 603 1385 637
rect 1419 603 1457 637
rect 1313 565 1491 603
rect 1347 531 1385 565
rect 1419 531 1457 565
rect 1313 493 1491 531
rect 1347 459 1385 493
rect 1419 459 1457 493
rect 1313 421 1491 459
rect 1347 387 1385 421
rect 1419 387 1457 421
rect 1313 349 1491 387
rect 1347 315 1385 349
rect 1419 315 1457 349
rect 1313 277 1491 315
rect 1347 243 1385 277
rect 1419 243 1457 277
rect 1313 205 1491 243
rect 1347 171 1385 205
rect 1419 171 1457 205
rect 1313 133 1491 171
rect 1347 99 1385 133
rect 1419 99 1457 133
rect 1313 83 1491 99
<< viali >>
rect 288 8132 322 8166
rect 360 8132 394 8166
rect 432 8132 466 8166
rect 504 8132 538 8166
rect 576 8132 610 8166
rect 648 8132 682 8166
rect 720 8132 754 8166
rect 792 8132 826 8166
rect 864 8132 898 8166
rect 936 8132 970 8166
rect 1008 8132 1042 8166
rect 74 8019 108 8053
rect 108 8019 146 8053
rect 146 8019 180 8053
rect 180 8019 218 8053
rect 218 8019 252 8053
rect 74 7981 252 8019
rect 74 7947 108 7981
rect 108 7947 146 7981
rect 146 7947 180 7981
rect 180 7947 218 7981
rect 218 7947 252 7981
rect 74 7909 252 7947
rect 74 7875 108 7909
rect 108 7875 146 7909
rect 146 7875 180 7909
rect 180 7875 218 7909
rect 218 7875 252 7909
rect 74 7837 252 7875
rect 74 7803 108 7837
rect 108 7803 146 7837
rect 146 7803 180 7837
rect 180 7803 218 7837
rect 218 7803 252 7837
rect 74 7765 252 7803
rect 74 7731 108 7765
rect 108 7731 146 7765
rect 146 7731 180 7765
rect 180 7731 218 7765
rect 218 7731 252 7765
rect 74 7693 252 7731
rect 74 7659 108 7693
rect 108 7659 146 7693
rect 146 7659 180 7693
rect 180 7659 218 7693
rect 218 7659 252 7693
rect 74 7621 252 7659
rect 74 7587 108 7621
rect 108 7587 146 7621
rect 146 7587 180 7621
rect 180 7587 218 7621
rect 218 7587 252 7621
rect 74 7549 252 7587
rect 74 7515 108 7549
rect 108 7515 146 7549
rect 146 7515 180 7549
rect 180 7515 218 7549
rect 218 7515 252 7549
rect 74 7477 252 7515
rect 74 7443 108 7477
rect 108 7443 146 7477
rect 146 7443 180 7477
rect 180 7443 218 7477
rect 218 7443 252 7477
rect 74 7405 252 7443
rect 74 7371 108 7405
rect 108 7371 146 7405
rect 146 7371 180 7405
rect 180 7371 218 7405
rect 218 7371 252 7405
rect 74 7333 252 7371
rect 74 7299 108 7333
rect 108 7299 146 7333
rect 146 7299 180 7333
rect 180 7299 218 7333
rect 218 7299 252 7333
rect 74 7261 252 7299
rect 74 7227 108 7261
rect 108 7227 146 7261
rect 146 7227 180 7261
rect 180 7227 218 7261
rect 218 7227 252 7261
rect 74 7189 252 7227
rect 74 7155 108 7189
rect 108 7155 146 7189
rect 146 7155 180 7189
rect 180 7155 218 7189
rect 218 7155 252 7189
rect 74 7117 252 7155
rect 74 7083 108 7117
rect 108 7083 146 7117
rect 146 7083 180 7117
rect 180 7083 218 7117
rect 218 7083 252 7117
rect 74 7045 252 7083
rect 74 7011 108 7045
rect 108 7011 146 7045
rect 146 7011 180 7045
rect 180 7011 218 7045
rect 218 7011 252 7045
rect 74 6973 252 7011
rect 74 6939 108 6973
rect 108 6939 146 6973
rect 146 6939 180 6973
rect 180 6939 218 6973
rect 218 6939 252 6973
rect 74 6901 252 6939
rect 74 6867 108 6901
rect 108 6867 146 6901
rect 146 6867 180 6901
rect 180 6867 218 6901
rect 218 6867 252 6901
rect 74 6829 252 6867
rect 74 6795 108 6829
rect 108 6795 146 6829
rect 146 6795 180 6829
rect 180 6795 218 6829
rect 218 6795 252 6829
rect 74 6757 252 6795
rect 74 6723 108 6757
rect 108 6723 146 6757
rect 146 6723 180 6757
rect 180 6723 218 6757
rect 218 6723 252 6757
rect 74 6685 252 6723
rect 74 6651 108 6685
rect 108 6651 146 6685
rect 146 6651 180 6685
rect 180 6651 218 6685
rect 218 6651 252 6685
rect 74 6613 252 6651
rect 74 6579 108 6613
rect 108 6579 146 6613
rect 146 6579 180 6613
rect 180 6579 218 6613
rect 218 6579 252 6613
rect 74 6541 252 6579
rect 74 6507 108 6541
rect 108 6507 146 6541
rect 146 6507 180 6541
rect 180 6507 218 6541
rect 218 6507 252 6541
rect 74 6469 252 6507
rect 74 6435 108 6469
rect 108 6435 146 6469
rect 146 6435 180 6469
rect 180 6435 218 6469
rect 218 6435 252 6469
rect 74 6397 252 6435
rect 74 6363 108 6397
rect 108 6363 146 6397
rect 146 6363 180 6397
rect 180 6363 218 6397
rect 218 6363 252 6397
rect 74 6325 252 6363
rect 74 6291 108 6325
rect 108 6291 146 6325
rect 146 6291 180 6325
rect 180 6291 218 6325
rect 218 6291 252 6325
rect 74 6253 252 6291
rect 74 6219 108 6253
rect 108 6219 146 6253
rect 146 6219 180 6253
rect 180 6219 218 6253
rect 218 6219 252 6253
rect 74 6181 252 6219
rect 74 6147 108 6181
rect 108 6147 146 6181
rect 146 6147 180 6181
rect 180 6147 218 6181
rect 218 6147 252 6181
rect 74 6109 252 6147
rect 74 6075 108 6109
rect 108 6075 146 6109
rect 146 6075 180 6109
rect 180 6075 218 6109
rect 218 6075 252 6109
rect 74 6037 252 6075
rect 74 6003 108 6037
rect 108 6003 146 6037
rect 146 6003 180 6037
rect 180 6003 218 6037
rect 218 6003 252 6037
rect 74 5965 252 6003
rect 74 5931 108 5965
rect 108 5931 146 5965
rect 146 5931 180 5965
rect 180 5931 218 5965
rect 218 5931 252 5965
rect 74 5893 252 5931
rect 74 5859 108 5893
rect 108 5859 146 5893
rect 146 5859 180 5893
rect 180 5859 218 5893
rect 218 5859 252 5893
rect 74 5821 252 5859
rect 74 5787 108 5821
rect 108 5787 146 5821
rect 146 5787 180 5821
rect 180 5787 218 5821
rect 218 5787 252 5821
rect 74 5749 252 5787
rect 74 5715 108 5749
rect 108 5715 146 5749
rect 146 5715 180 5749
rect 180 5715 218 5749
rect 218 5715 252 5749
rect 74 5677 252 5715
rect 74 5643 108 5677
rect 108 5643 146 5677
rect 146 5643 180 5677
rect 180 5643 218 5677
rect 218 5643 252 5677
rect 74 5605 252 5643
rect 74 5571 108 5605
rect 108 5571 146 5605
rect 146 5571 180 5605
rect 180 5571 218 5605
rect 218 5571 252 5605
rect 74 5533 252 5571
rect 74 5499 108 5533
rect 108 5499 146 5533
rect 146 5499 180 5533
rect 180 5499 218 5533
rect 218 5499 252 5533
rect 74 5461 252 5499
rect 74 5427 108 5461
rect 108 5427 146 5461
rect 146 5427 180 5461
rect 180 5427 218 5461
rect 218 5427 252 5461
rect 74 5389 252 5427
rect 74 5355 108 5389
rect 108 5355 146 5389
rect 146 5355 180 5389
rect 180 5355 218 5389
rect 218 5355 252 5389
rect 74 5317 252 5355
rect 74 5283 108 5317
rect 108 5283 146 5317
rect 146 5283 180 5317
rect 180 5283 218 5317
rect 218 5283 252 5317
rect 74 5245 252 5283
rect 74 5211 108 5245
rect 108 5211 146 5245
rect 146 5211 180 5245
rect 180 5211 218 5245
rect 218 5211 252 5245
rect 74 5173 252 5211
rect 74 5139 108 5173
rect 108 5139 146 5173
rect 146 5139 180 5173
rect 180 5139 218 5173
rect 218 5139 252 5173
rect 74 5101 252 5139
rect 74 5067 108 5101
rect 108 5067 146 5101
rect 146 5067 180 5101
rect 180 5067 218 5101
rect 218 5067 252 5101
rect 74 5029 252 5067
rect 74 4995 108 5029
rect 108 4995 146 5029
rect 146 4995 180 5029
rect 180 4995 218 5029
rect 218 4995 252 5029
rect 74 4957 252 4995
rect 74 4923 108 4957
rect 108 4923 146 4957
rect 146 4923 180 4957
rect 180 4923 218 4957
rect 218 4923 252 4957
rect 74 4885 252 4923
rect 74 4851 108 4885
rect 108 4851 146 4885
rect 146 4851 180 4885
rect 180 4851 218 4885
rect 218 4851 252 4885
rect 74 4813 252 4851
rect 74 4779 108 4813
rect 108 4779 146 4813
rect 146 4779 180 4813
rect 180 4779 218 4813
rect 218 4779 252 4813
rect 74 4741 252 4779
rect 74 4707 108 4741
rect 108 4707 146 4741
rect 146 4707 180 4741
rect 180 4707 218 4741
rect 218 4707 252 4741
rect 74 4669 252 4707
rect 74 4635 108 4669
rect 108 4635 146 4669
rect 146 4635 180 4669
rect 180 4635 218 4669
rect 218 4635 252 4669
rect 74 4597 252 4635
rect 74 4563 108 4597
rect 108 4563 146 4597
rect 146 4563 180 4597
rect 180 4563 218 4597
rect 218 4563 252 4597
rect 74 4525 252 4563
rect 74 4491 108 4525
rect 108 4491 146 4525
rect 146 4491 180 4525
rect 180 4491 218 4525
rect 218 4491 252 4525
rect 74 4453 252 4491
rect 74 4419 108 4453
rect 108 4419 146 4453
rect 146 4419 180 4453
rect 180 4419 218 4453
rect 218 4419 252 4453
rect 74 4381 252 4419
rect 74 4347 108 4381
rect 108 4347 146 4381
rect 146 4347 180 4381
rect 180 4347 218 4381
rect 218 4347 252 4381
rect 74 4309 252 4347
rect 74 4275 108 4309
rect 108 4275 146 4309
rect 146 4275 180 4309
rect 180 4275 218 4309
rect 218 4275 252 4309
rect 74 4237 252 4275
rect 74 4203 108 4237
rect 108 4203 146 4237
rect 146 4203 180 4237
rect 180 4203 218 4237
rect 218 4203 252 4237
rect 74 4165 252 4203
rect 74 4131 108 4165
rect 108 4131 146 4165
rect 146 4131 180 4165
rect 180 4131 218 4165
rect 218 4131 252 4165
rect 74 4093 252 4131
rect 74 4059 108 4093
rect 108 4059 146 4093
rect 146 4059 180 4093
rect 180 4059 218 4093
rect 218 4059 252 4093
rect 74 4021 252 4059
rect 74 3987 108 4021
rect 108 3987 146 4021
rect 146 3987 180 4021
rect 180 3987 218 4021
rect 218 3987 252 4021
rect 74 3949 252 3987
rect 74 3915 108 3949
rect 108 3915 146 3949
rect 146 3915 180 3949
rect 180 3915 218 3949
rect 218 3915 252 3949
rect 74 3877 252 3915
rect 74 3843 108 3877
rect 108 3843 146 3877
rect 146 3843 180 3877
rect 180 3843 218 3877
rect 218 3843 252 3877
rect 74 3805 252 3843
rect 74 3771 108 3805
rect 108 3771 146 3805
rect 146 3771 180 3805
rect 180 3771 218 3805
rect 218 3771 252 3805
rect 74 3733 252 3771
rect 74 3699 108 3733
rect 108 3699 146 3733
rect 146 3699 180 3733
rect 180 3699 218 3733
rect 218 3699 252 3733
rect 74 3661 252 3699
rect 74 3627 108 3661
rect 108 3627 146 3661
rect 146 3627 180 3661
rect 180 3627 218 3661
rect 218 3627 252 3661
rect 74 3589 252 3627
rect 74 3555 108 3589
rect 108 3555 146 3589
rect 146 3555 180 3589
rect 180 3555 218 3589
rect 218 3555 252 3589
rect 74 3517 252 3555
rect 74 3483 108 3517
rect 108 3483 146 3517
rect 146 3483 180 3517
rect 180 3483 218 3517
rect 218 3483 252 3517
rect 74 3445 252 3483
rect 74 3411 108 3445
rect 108 3411 146 3445
rect 146 3411 180 3445
rect 180 3411 218 3445
rect 218 3411 252 3445
rect 74 3373 252 3411
rect 74 3339 108 3373
rect 108 3339 146 3373
rect 146 3339 180 3373
rect 180 3339 218 3373
rect 218 3339 252 3373
rect 74 3301 252 3339
rect 74 3267 108 3301
rect 108 3267 146 3301
rect 146 3267 180 3301
rect 180 3267 218 3301
rect 218 3267 252 3301
rect 74 3229 252 3267
rect 74 3195 108 3229
rect 108 3195 146 3229
rect 146 3195 180 3229
rect 180 3195 218 3229
rect 218 3195 252 3229
rect 74 3157 252 3195
rect 74 3123 108 3157
rect 108 3123 146 3157
rect 146 3123 180 3157
rect 180 3123 218 3157
rect 218 3123 252 3157
rect 74 3085 252 3123
rect 74 3051 108 3085
rect 108 3051 146 3085
rect 146 3051 180 3085
rect 180 3051 218 3085
rect 218 3051 252 3085
rect 74 3013 252 3051
rect 74 2979 108 3013
rect 108 2979 146 3013
rect 146 2979 180 3013
rect 180 2979 218 3013
rect 218 2979 252 3013
rect 74 2941 252 2979
rect 74 2907 108 2941
rect 108 2907 146 2941
rect 146 2907 180 2941
rect 180 2907 218 2941
rect 218 2907 252 2941
rect 74 2869 252 2907
rect 74 2835 108 2869
rect 108 2835 146 2869
rect 146 2835 180 2869
rect 180 2835 218 2869
rect 218 2835 252 2869
rect 74 2797 252 2835
rect 74 2763 108 2797
rect 108 2763 146 2797
rect 146 2763 180 2797
rect 180 2763 218 2797
rect 218 2763 252 2797
rect 74 2725 252 2763
rect 74 2691 108 2725
rect 108 2691 146 2725
rect 146 2691 180 2725
rect 180 2691 218 2725
rect 218 2691 252 2725
rect 74 2653 252 2691
rect 74 2619 108 2653
rect 108 2619 146 2653
rect 146 2619 180 2653
rect 180 2619 218 2653
rect 218 2619 252 2653
rect 74 2581 252 2619
rect 74 2547 108 2581
rect 108 2547 146 2581
rect 146 2547 180 2581
rect 180 2547 218 2581
rect 218 2547 252 2581
rect 74 2509 252 2547
rect 74 2475 108 2509
rect 108 2475 146 2509
rect 146 2475 180 2509
rect 180 2475 218 2509
rect 218 2475 252 2509
rect 74 2437 252 2475
rect 74 2403 108 2437
rect 108 2403 146 2437
rect 146 2403 180 2437
rect 180 2403 218 2437
rect 218 2403 252 2437
rect 74 2365 252 2403
rect 74 2331 108 2365
rect 108 2331 146 2365
rect 146 2331 180 2365
rect 180 2331 218 2365
rect 218 2331 252 2365
rect 74 2293 252 2331
rect 74 2259 108 2293
rect 108 2259 146 2293
rect 146 2259 180 2293
rect 180 2259 218 2293
rect 218 2259 252 2293
rect 74 2221 252 2259
rect 74 2187 108 2221
rect 108 2187 146 2221
rect 146 2187 180 2221
rect 180 2187 218 2221
rect 218 2187 252 2221
rect 74 2149 252 2187
rect 74 2115 108 2149
rect 108 2115 146 2149
rect 146 2115 180 2149
rect 180 2115 218 2149
rect 218 2115 252 2149
rect 74 2077 252 2115
rect 74 2043 108 2077
rect 108 2043 146 2077
rect 146 2043 180 2077
rect 180 2043 218 2077
rect 218 2043 252 2077
rect 74 2005 252 2043
rect 74 1971 108 2005
rect 108 1971 146 2005
rect 146 1971 180 2005
rect 180 1971 218 2005
rect 218 1971 252 2005
rect 74 1933 252 1971
rect 74 1899 108 1933
rect 108 1899 146 1933
rect 146 1899 180 1933
rect 180 1899 218 1933
rect 218 1899 252 1933
rect 74 1861 252 1899
rect 74 1827 108 1861
rect 108 1827 146 1861
rect 146 1827 180 1861
rect 180 1827 218 1861
rect 218 1827 252 1861
rect 74 1789 252 1827
rect 74 1755 108 1789
rect 108 1755 146 1789
rect 146 1755 180 1789
rect 180 1755 218 1789
rect 218 1755 252 1789
rect 74 1717 252 1755
rect 74 1683 108 1717
rect 108 1683 146 1717
rect 146 1683 180 1717
rect 180 1683 218 1717
rect 218 1683 252 1717
rect 74 1645 252 1683
rect 74 1611 108 1645
rect 108 1611 146 1645
rect 146 1611 180 1645
rect 180 1611 218 1645
rect 218 1611 252 1645
rect 74 1573 252 1611
rect 74 1539 108 1573
rect 108 1539 146 1573
rect 146 1539 180 1573
rect 180 1539 218 1573
rect 218 1539 252 1573
rect 74 1501 252 1539
rect 74 1467 108 1501
rect 108 1467 146 1501
rect 146 1467 180 1501
rect 180 1467 218 1501
rect 218 1467 252 1501
rect 74 1429 252 1467
rect 74 1395 108 1429
rect 108 1395 146 1429
rect 146 1395 180 1429
rect 180 1395 218 1429
rect 218 1395 252 1429
rect 74 1357 252 1395
rect 74 1323 108 1357
rect 108 1323 146 1357
rect 146 1323 180 1357
rect 180 1323 218 1357
rect 218 1323 252 1357
rect 74 1285 252 1323
rect 74 1251 108 1285
rect 108 1251 146 1285
rect 146 1251 180 1285
rect 180 1251 218 1285
rect 218 1251 252 1285
rect 74 1213 252 1251
rect 74 1179 108 1213
rect 108 1179 146 1213
rect 146 1179 180 1213
rect 180 1179 218 1213
rect 218 1179 252 1213
rect 74 1141 252 1179
rect 74 1107 108 1141
rect 108 1107 146 1141
rect 146 1107 180 1141
rect 180 1107 218 1141
rect 218 1107 252 1141
rect 74 1069 252 1107
rect 74 1035 108 1069
rect 108 1035 146 1069
rect 146 1035 180 1069
rect 180 1035 218 1069
rect 218 1035 252 1069
rect 74 997 252 1035
rect 74 963 108 997
rect 108 963 146 997
rect 146 963 180 997
rect 180 963 218 997
rect 218 963 252 997
rect 74 925 252 963
rect 74 891 108 925
rect 108 891 146 925
rect 146 891 180 925
rect 180 891 218 925
rect 218 891 252 925
rect 74 853 252 891
rect 74 819 108 853
rect 108 819 146 853
rect 146 819 180 853
rect 180 819 218 853
rect 218 819 252 853
rect 74 781 252 819
rect 74 747 108 781
rect 108 747 146 781
rect 146 747 180 781
rect 180 747 218 781
rect 218 747 252 781
rect 74 709 252 747
rect 74 675 108 709
rect 108 675 146 709
rect 146 675 180 709
rect 180 675 218 709
rect 218 675 252 709
rect 74 637 252 675
rect 74 603 108 637
rect 108 603 146 637
rect 146 603 180 637
rect 180 603 218 637
rect 218 603 252 637
rect 74 565 252 603
rect 74 531 108 565
rect 108 531 146 565
rect 146 531 180 565
rect 180 531 218 565
rect 218 531 252 565
rect 74 493 252 531
rect 74 459 108 493
rect 108 459 146 493
rect 146 459 180 493
rect 180 459 218 493
rect 218 459 252 493
rect 74 421 252 459
rect 74 387 108 421
rect 108 387 146 421
rect 146 387 180 421
rect 180 387 218 421
rect 218 387 252 421
rect 74 349 252 387
rect 74 315 108 349
rect 108 315 146 349
rect 146 315 180 349
rect 180 315 218 349
rect 218 315 252 349
rect 74 277 252 315
rect 74 243 108 277
rect 108 243 146 277
rect 146 243 180 277
rect 180 243 218 277
rect 218 243 252 277
rect 74 205 252 243
rect 74 171 108 205
rect 108 171 146 205
rect 146 171 180 205
rect 180 171 218 205
rect 218 171 252 205
rect 74 133 252 171
rect 74 99 108 133
rect 108 99 146 133
rect 146 99 180 133
rect 180 99 218 133
rect 218 99 252 133
rect 1078 8019 1112 8053
rect 1112 8019 1150 8053
rect 1150 8019 1184 8053
rect 1184 8019 1222 8053
rect 1222 8019 1256 8053
rect 1078 7981 1256 8019
rect 1078 7947 1112 7981
rect 1112 7947 1150 7981
rect 1150 7947 1184 7981
rect 1184 7947 1222 7981
rect 1222 7947 1256 7981
rect 1078 7909 1256 7947
rect 1078 7875 1112 7909
rect 1112 7875 1150 7909
rect 1150 7875 1184 7909
rect 1184 7875 1222 7909
rect 1222 7875 1256 7909
rect 1078 7837 1256 7875
rect 1078 7803 1112 7837
rect 1112 7803 1150 7837
rect 1150 7803 1184 7837
rect 1184 7803 1222 7837
rect 1222 7803 1256 7837
rect 1078 7765 1256 7803
rect 1078 7731 1112 7765
rect 1112 7731 1150 7765
rect 1150 7731 1184 7765
rect 1184 7731 1222 7765
rect 1222 7731 1256 7765
rect 1078 7693 1256 7731
rect 1078 7659 1112 7693
rect 1112 7659 1150 7693
rect 1150 7659 1184 7693
rect 1184 7659 1222 7693
rect 1222 7659 1256 7693
rect 1078 7621 1256 7659
rect 1078 7587 1112 7621
rect 1112 7587 1150 7621
rect 1150 7587 1184 7621
rect 1184 7587 1222 7621
rect 1222 7587 1256 7621
rect 1078 7549 1256 7587
rect 1078 7515 1112 7549
rect 1112 7515 1150 7549
rect 1150 7515 1184 7549
rect 1184 7515 1222 7549
rect 1222 7515 1256 7549
rect 1078 7477 1256 7515
rect 1078 7443 1112 7477
rect 1112 7443 1150 7477
rect 1150 7443 1184 7477
rect 1184 7443 1222 7477
rect 1222 7443 1256 7477
rect 1078 7405 1256 7443
rect 1078 7371 1112 7405
rect 1112 7371 1150 7405
rect 1150 7371 1184 7405
rect 1184 7371 1222 7405
rect 1222 7371 1256 7405
rect 1078 7333 1256 7371
rect 1078 7299 1112 7333
rect 1112 7299 1150 7333
rect 1150 7299 1184 7333
rect 1184 7299 1222 7333
rect 1222 7299 1256 7333
rect 1078 7261 1256 7299
rect 1078 7227 1112 7261
rect 1112 7227 1150 7261
rect 1150 7227 1184 7261
rect 1184 7227 1222 7261
rect 1222 7227 1256 7261
rect 1078 7189 1256 7227
rect 1078 7155 1112 7189
rect 1112 7155 1150 7189
rect 1150 7155 1184 7189
rect 1184 7155 1222 7189
rect 1222 7155 1256 7189
rect 1078 7117 1256 7155
rect 1078 7083 1112 7117
rect 1112 7083 1150 7117
rect 1150 7083 1184 7117
rect 1184 7083 1222 7117
rect 1222 7083 1256 7117
rect 1078 7045 1256 7083
rect 1078 7011 1112 7045
rect 1112 7011 1150 7045
rect 1150 7011 1184 7045
rect 1184 7011 1222 7045
rect 1222 7011 1256 7045
rect 1078 6973 1256 7011
rect 1078 6939 1112 6973
rect 1112 6939 1150 6973
rect 1150 6939 1184 6973
rect 1184 6939 1222 6973
rect 1222 6939 1256 6973
rect 1078 6901 1256 6939
rect 1078 6867 1112 6901
rect 1112 6867 1150 6901
rect 1150 6867 1184 6901
rect 1184 6867 1222 6901
rect 1222 6867 1256 6901
rect 1078 6829 1256 6867
rect 1078 6795 1112 6829
rect 1112 6795 1150 6829
rect 1150 6795 1184 6829
rect 1184 6795 1222 6829
rect 1222 6795 1256 6829
rect 1078 6757 1256 6795
rect 1078 6723 1112 6757
rect 1112 6723 1150 6757
rect 1150 6723 1184 6757
rect 1184 6723 1222 6757
rect 1222 6723 1256 6757
rect 1078 6685 1256 6723
rect 1078 6651 1112 6685
rect 1112 6651 1150 6685
rect 1150 6651 1184 6685
rect 1184 6651 1222 6685
rect 1222 6651 1256 6685
rect 1078 6613 1256 6651
rect 1078 6579 1112 6613
rect 1112 6579 1150 6613
rect 1150 6579 1184 6613
rect 1184 6579 1222 6613
rect 1222 6579 1256 6613
rect 1078 6541 1256 6579
rect 1078 6507 1112 6541
rect 1112 6507 1150 6541
rect 1150 6507 1184 6541
rect 1184 6507 1222 6541
rect 1222 6507 1256 6541
rect 1078 6469 1256 6507
rect 1078 6435 1112 6469
rect 1112 6435 1150 6469
rect 1150 6435 1184 6469
rect 1184 6435 1222 6469
rect 1222 6435 1256 6469
rect 1078 6397 1256 6435
rect 1078 6363 1112 6397
rect 1112 6363 1150 6397
rect 1150 6363 1184 6397
rect 1184 6363 1222 6397
rect 1222 6363 1256 6397
rect 1078 6325 1256 6363
rect 1078 6291 1112 6325
rect 1112 6291 1150 6325
rect 1150 6291 1184 6325
rect 1184 6291 1222 6325
rect 1222 6291 1256 6325
rect 1078 6253 1256 6291
rect 1078 6219 1112 6253
rect 1112 6219 1150 6253
rect 1150 6219 1184 6253
rect 1184 6219 1222 6253
rect 1222 6219 1256 6253
rect 1078 6181 1256 6219
rect 1078 6147 1112 6181
rect 1112 6147 1150 6181
rect 1150 6147 1184 6181
rect 1184 6147 1222 6181
rect 1222 6147 1256 6181
rect 1078 6109 1256 6147
rect 1078 6075 1112 6109
rect 1112 6075 1150 6109
rect 1150 6075 1184 6109
rect 1184 6075 1222 6109
rect 1222 6075 1256 6109
rect 1078 6037 1256 6075
rect 1078 6003 1112 6037
rect 1112 6003 1150 6037
rect 1150 6003 1184 6037
rect 1184 6003 1222 6037
rect 1222 6003 1256 6037
rect 1078 5965 1256 6003
rect 1078 5931 1112 5965
rect 1112 5931 1150 5965
rect 1150 5931 1184 5965
rect 1184 5931 1222 5965
rect 1222 5931 1256 5965
rect 1078 5893 1256 5931
rect 1078 5859 1112 5893
rect 1112 5859 1150 5893
rect 1150 5859 1184 5893
rect 1184 5859 1222 5893
rect 1222 5859 1256 5893
rect 1078 5821 1256 5859
rect 1078 5787 1112 5821
rect 1112 5787 1150 5821
rect 1150 5787 1184 5821
rect 1184 5787 1222 5821
rect 1222 5787 1256 5821
rect 1078 5749 1256 5787
rect 1078 5715 1112 5749
rect 1112 5715 1150 5749
rect 1150 5715 1184 5749
rect 1184 5715 1222 5749
rect 1222 5715 1256 5749
rect 1078 5677 1256 5715
rect 1078 5643 1112 5677
rect 1112 5643 1150 5677
rect 1150 5643 1184 5677
rect 1184 5643 1222 5677
rect 1222 5643 1256 5677
rect 1078 5605 1256 5643
rect 1078 5571 1112 5605
rect 1112 5571 1150 5605
rect 1150 5571 1184 5605
rect 1184 5571 1222 5605
rect 1222 5571 1256 5605
rect 1078 5533 1256 5571
rect 1078 5499 1112 5533
rect 1112 5499 1150 5533
rect 1150 5499 1184 5533
rect 1184 5499 1222 5533
rect 1222 5499 1256 5533
rect 1078 5461 1256 5499
rect 1078 5427 1112 5461
rect 1112 5427 1150 5461
rect 1150 5427 1184 5461
rect 1184 5427 1222 5461
rect 1222 5427 1256 5461
rect 1078 5389 1256 5427
rect 1078 5355 1112 5389
rect 1112 5355 1150 5389
rect 1150 5355 1184 5389
rect 1184 5355 1222 5389
rect 1222 5355 1256 5389
rect 1078 5317 1256 5355
rect 1078 5283 1112 5317
rect 1112 5283 1150 5317
rect 1150 5283 1184 5317
rect 1184 5283 1222 5317
rect 1222 5283 1256 5317
rect 1078 5245 1256 5283
rect 1078 5211 1112 5245
rect 1112 5211 1150 5245
rect 1150 5211 1184 5245
rect 1184 5211 1222 5245
rect 1222 5211 1256 5245
rect 1078 5173 1256 5211
rect 1078 5139 1112 5173
rect 1112 5139 1150 5173
rect 1150 5139 1184 5173
rect 1184 5139 1222 5173
rect 1222 5139 1256 5173
rect 1078 5101 1256 5139
rect 1078 5067 1112 5101
rect 1112 5067 1150 5101
rect 1150 5067 1184 5101
rect 1184 5067 1222 5101
rect 1222 5067 1256 5101
rect 1078 5029 1256 5067
rect 1078 4995 1112 5029
rect 1112 4995 1150 5029
rect 1150 4995 1184 5029
rect 1184 4995 1222 5029
rect 1222 4995 1256 5029
rect 1078 4957 1256 4995
rect 1078 4923 1112 4957
rect 1112 4923 1150 4957
rect 1150 4923 1184 4957
rect 1184 4923 1222 4957
rect 1222 4923 1256 4957
rect 1078 4885 1256 4923
rect 1078 4851 1112 4885
rect 1112 4851 1150 4885
rect 1150 4851 1184 4885
rect 1184 4851 1222 4885
rect 1222 4851 1256 4885
rect 1078 4813 1256 4851
rect 1078 4779 1112 4813
rect 1112 4779 1150 4813
rect 1150 4779 1184 4813
rect 1184 4779 1222 4813
rect 1222 4779 1256 4813
rect 1078 4741 1256 4779
rect 1078 4707 1112 4741
rect 1112 4707 1150 4741
rect 1150 4707 1184 4741
rect 1184 4707 1222 4741
rect 1222 4707 1256 4741
rect 1078 4669 1256 4707
rect 1078 4635 1112 4669
rect 1112 4635 1150 4669
rect 1150 4635 1184 4669
rect 1184 4635 1222 4669
rect 1222 4635 1256 4669
rect 1078 4597 1256 4635
rect 1078 4563 1112 4597
rect 1112 4563 1150 4597
rect 1150 4563 1184 4597
rect 1184 4563 1222 4597
rect 1222 4563 1256 4597
rect 1078 4525 1256 4563
rect 1078 4491 1112 4525
rect 1112 4491 1150 4525
rect 1150 4491 1184 4525
rect 1184 4491 1222 4525
rect 1222 4491 1256 4525
rect 1078 4453 1256 4491
rect 1078 4419 1112 4453
rect 1112 4419 1150 4453
rect 1150 4419 1184 4453
rect 1184 4419 1222 4453
rect 1222 4419 1256 4453
rect 1078 4381 1256 4419
rect 1078 4347 1112 4381
rect 1112 4347 1150 4381
rect 1150 4347 1184 4381
rect 1184 4347 1222 4381
rect 1222 4347 1256 4381
rect 1078 4309 1256 4347
rect 1078 4275 1112 4309
rect 1112 4275 1150 4309
rect 1150 4275 1184 4309
rect 1184 4275 1222 4309
rect 1222 4275 1256 4309
rect 1078 4237 1256 4275
rect 1078 4203 1112 4237
rect 1112 4203 1150 4237
rect 1150 4203 1184 4237
rect 1184 4203 1222 4237
rect 1222 4203 1256 4237
rect 1078 4165 1256 4203
rect 1078 4131 1112 4165
rect 1112 4131 1150 4165
rect 1150 4131 1184 4165
rect 1184 4131 1222 4165
rect 1222 4131 1256 4165
rect 1078 4093 1256 4131
rect 1078 4059 1112 4093
rect 1112 4059 1150 4093
rect 1150 4059 1184 4093
rect 1184 4059 1222 4093
rect 1222 4059 1256 4093
rect 1078 4021 1256 4059
rect 1078 3987 1112 4021
rect 1112 3987 1150 4021
rect 1150 3987 1184 4021
rect 1184 3987 1222 4021
rect 1222 3987 1256 4021
rect 1078 3949 1256 3987
rect 1078 3915 1112 3949
rect 1112 3915 1150 3949
rect 1150 3915 1184 3949
rect 1184 3915 1222 3949
rect 1222 3915 1256 3949
rect 1078 3877 1256 3915
rect 1078 3843 1112 3877
rect 1112 3843 1150 3877
rect 1150 3843 1184 3877
rect 1184 3843 1222 3877
rect 1222 3843 1256 3877
rect 1078 3805 1256 3843
rect 1078 3771 1112 3805
rect 1112 3771 1150 3805
rect 1150 3771 1184 3805
rect 1184 3771 1222 3805
rect 1222 3771 1256 3805
rect 1078 3733 1256 3771
rect 1078 3699 1112 3733
rect 1112 3699 1150 3733
rect 1150 3699 1184 3733
rect 1184 3699 1222 3733
rect 1222 3699 1256 3733
rect 1078 3661 1256 3699
rect 1078 3627 1112 3661
rect 1112 3627 1150 3661
rect 1150 3627 1184 3661
rect 1184 3627 1222 3661
rect 1222 3627 1256 3661
rect 1078 3589 1256 3627
rect 1078 3555 1112 3589
rect 1112 3555 1150 3589
rect 1150 3555 1184 3589
rect 1184 3555 1222 3589
rect 1222 3555 1256 3589
rect 1078 3517 1256 3555
rect 1078 3483 1112 3517
rect 1112 3483 1150 3517
rect 1150 3483 1184 3517
rect 1184 3483 1222 3517
rect 1222 3483 1256 3517
rect 1078 3445 1256 3483
rect 1078 3411 1112 3445
rect 1112 3411 1150 3445
rect 1150 3411 1184 3445
rect 1184 3411 1222 3445
rect 1222 3411 1256 3445
rect 1078 3373 1256 3411
rect 1078 3339 1112 3373
rect 1112 3339 1150 3373
rect 1150 3339 1184 3373
rect 1184 3339 1222 3373
rect 1222 3339 1256 3373
rect 1078 3301 1256 3339
rect 1078 3267 1112 3301
rect 1112 3267 1150 3301
rect 1150 3267 1184 3301
rect 1184 3267 1222 3301
rect 1222 3267 1256 3301
rect 1078 3229 1256 3267
rect 1078 3195 1112 3229
rect 1112 3195 1150 3229
rect 1150 3195 1184 3229
rect 1184 3195 1222 3229
rect 1222 3195 1256 3229
rect 1078 3157 1256 3195
rect 1078 3123 1112 3157
rect 1112 3123 1150 3157
rect 1150 3123 1184 3157
rect 1184 3123 1222 3157
rect 1222 3123 1256 3157
rect 1078 3085 1256 3123
rect 1078 3051 1112 3085
rect 1112 3051 1150 3085
rect 1150 3051 1184 3085
rect 1184 3051 1222 3085
rect 1222 3051 1256 3085
rect 1078 3013 1256 3051
rect 1078 2979 1112 3013
rect 1112 2979 1150 3013
rect 1150 2979 1184 3013
rect 1184 2979 1222 3013
rect 1222 2979 1256 3013
rect 1078 2941 1256 2979
rect 1078 2907 1112 2941
rect 1112 2907 1150 2941
rect 1150 2907 1184 2941
rect 1184 2907 1222 2941
rect 1222 2907 1256 2941
rect 1078 2869 1256 2907
rect 1078 2835 1112 2869
rect 1112 2835 1150 2869
rect 1150 2835 1184 2869
rect 1184 2835 1222 2869
rect 1222 2835 1256 2869
rect 1078 2797 1256 2835
rect 1078 2763 1112 2797
rect 1112 2763 1150 2797
rect 1150 2763 1184 2797
rect 1184 2763 1222 2797
rect 1222 2763 1256 2797
rect 1078 2725 1256 2763
rect 1078 2691 1112 2725
rect 1112 2691 1150 2725
rect 1150 2691 1184 2725
rect 1184 2691 1222 2725
rect 1222 2691 1256 2725
rect 1078 2653 1256 2691
rect 1078 2619 1112 2653
rect 1112 2619 1150 2653
rect 1150 2619 1184 2653
rect 1184 2619 1222 2653
rect 1222 2619 1256 2653
rect 1078 2581 1256 2619
rect 1078 2547 1112 2581
rect 1112 2547 1150 2581
rect 1150 2547 1184 2581
rect 1184 2547 1222 2581
rect 1222 2547 1256 2581
rect 1078 2509 1256 2547
rect 1078 2475 1112 2509
rect 1112 2475 1150 2509
rect 1150 2475 1184 2509
rect 1184 2475 1222 2509
rect 1222 2475 1256 2509
rect 1078 2437 1256 2475
rect 1078 2403 1112 2437
rect 1112 2403 1150 2437
rect 1150 2403 1184 2437
rect 1184 2403 1222 2437
rect 1222 2403 1256 2437
rect 1078 2365 1256 2403
rect 1078 2331 1112 2365
rect 1112 2331 1150 2365
rect 1150 2331 1184 2365
rect 1184 2331 1222 2365
rect 1222 2331 1256 2365
rect 1078 2293 1256 2331
rect 1078 2259 1112 2293
rect 1112 2259 1150 2293
rect 1150 2259 1184 2293
rect 1184 2259 1222 2293
rect 1222 2259 1256 2293
rect 1078 2221 1256 2259
rect 1078 2187 1112 2221
rect 1112 2187 1150 2221
rect 1150 2187 1184 2221
rect 1184 2187 1222 2221
rect 1222 2187 1256 2221
rect 1078 2149 1256 2187
rect 1078 2115 1112 2149
rect 1112 2115 1150 2149
rect 1150 2115 1184 2149
rect 1184 2115 1222 2149
rect 1222 2115 1256 2149
rect 1078 2077 1256 2115
rect 1078 2043 1112 2077
rect 1112 2043 1150 2077
rect 1150 2043 1184 2077
rect 1184 2043 1222 2077
rect 1222 2043 1256 2077
rect 1078 2005 1256 2043
rect 1078 1971 1112 2005
rect 1112 1971 1150 2005
rect 1150 1971 1184 2005
rect 1184 1971 1222 2005
rect 1222 1971 1256 2005
rect 1078 1933 1256 1971
rect 1078 1899 1112 1933
rect 1112 1899 1150 1933
rect 1150 1899 1184 1933
rect 1184 1899 1222 1933
rect 1222 1899 1256 1933
rect 1078 1861 1256 1899
rect 1078 1827 1112 1861
rect 1112 1827 1150 1861
rect 1150 1827 1184 1861
rect 1184 1827 1222 1861
rect 1222 1827 1256 1861
rect 1078 1789 1256 1827
rect 1078 1755 1112 1789
rect 1112 1755 1150 1789
rect 1150 1755 1184 1789
rect 1184 1755 1222 1789
rect 1222 1755 1256 1789
rect 1078 1717 1256 1755
rect 1078 1683 1112 1717
rect 1112 1683 1150 1717
rect 1150 1683 1184 1717
rect 1184 1683 1222 1717
rect 1222 1683 1256 1717
rect 1078 1645 1256 1683
rect 1078 1611 1112 1645
rect 1112 1611 1150 1645
rect 1150 1611 1184 1645
rect 1184 1611 1222 1645
rect 1222 1611 1256 1645
rect 1078 1573 1256 1611
rect 1078 1539 1112 1573
rect 1112 1539 1150 1573
rect 1150 1539 1184 1573
rect 1184 1539 1222 1573
rect 1222 1539 1256 1573
rect 1078 1501 1256 1539
rect 1078 1467 1112 1501
rect 1112 1467 1150 1501
rect 1150 1467 1184 1501
rect 1184 1467 1222 1501
rect 1222 1467 1256 1501
rect 1078 1429 1256 1467
rect 1078 1395 1112 1429
rect 1112 1395 1150 1429
rect 1150 1395 1184 1429
rect 1184 1395 1222 1429
rect 1222 1395 1256 1429
rect 1078 1357 1256 1395
rect 1078 1323 1112 1357
rect 1112 1323 1150 1357
rect 1150 1323 1184 1357
rect 1184 1323 1222 1357
rect 1222 1323 1256 1357
rect 1078 1285 1256 1323
rect 1078 1251 1112 1285
rect 1112 1251 1150 1285
rect 1150 1251 1184 1285
rect 1184 1251 1222 1285
rect 1222 1251 1256 1285
rect 1078 1213 1256 1251
rect 1078 1179 1112 1213
rect 1112 1179 1150 1213
rect 1150 1179 1184 1213
rect 1184 1179 1222 1213
rect 1222 1179 1256 1213
rect 1078 1141 1256 1179
rect 1078 1107 1112 1141
rect 1112 1107 1150 1141
rect 1150 1107 1184 1141
rect 1184 1107 1222 1141
rect 1222 1107 1256 1141
rect 1078 1069 1256 1107
rect 1078 1035 1112 1069
rect 1112 1035 1150 1069
rect 1150 1035 1184 1069
rect 1184 1035 1222 1069
rect 1222 1035 1256 1069
rect 1078 997 1256 1035
rect 1078 963 1112 997
rect 1112 963 1150 997
rect 1150 963 1184 997
rect 1184 963 1222 997
rect 1222 963 1256 997
rect 1078 925 1256 963
rect 1078 891 1112 925
rect 1112 891 1150 925
rect 1150 891 1184 925
rect 1184 891 1222 925
rect 1222 891 1256 925
rect 1078 853 1256 891
rect 1078 819 1112 853
rect 1112 819 1150 853
rect 1150 819 1184 853
rect 1184 819 1222 853
rect 1222 819 1256 853
rect 1078 781 1256 819
rect 1078 747 1112 781
rect 1112 747 1150 781
rect 1150 747 1184 781
rect 1184 747 1222 781
rect 1222 747 1256 781
rect 1078 709 1256 747
rect 1078 675 1112 709
rect 1112 675 1150 709
rect 1150 675 1184 709
rect 1184 675 1222 709
rect 1222 675 1256 709
rect 1078 637 1256 675
rect 1078 603 1112 637
rect 1112 603 1150 637
rect 1150 603 1184 637
rect 1184 603 1222 637
rect 1222 603 1256 637
rect 1078 565 1256 603
rect 1078 531 1112 565
rect 1112 531 1150 565
rect 1150 531 1184 565
rect 1184 531 1222 565
rect 1222 531 1256 565
rect 1078 493 1256 531
rect 1078 459 1112 493
rect 1112 459 1150 493
rect 1150 459 1184 493
rect 1184 459 1222 493
rect 1222 459 1256 493
rect 1078 421 1256 459
rect 1078 387 1112 421
rect 1112 387 1150 421
rect 1150 387 1184 421
rect 1184 387 1222 421
rect 1222 387 1256 421
rect 1078 349 1256 387
rect 1078 315 1112 349
rect 1112 315 1150 349
rect 1150 315 1184 349
rect 1184 315 1222 349
rect 1222 315 1256 349
rect 1078 277 1256 315
rect 1078 243 1112 277
rect 1112 243 1150 277
rect 1150 243 1184 277
rect 1184 243 1222 277
rect 1222 243 1256 277
rect 1078 205 1256 243
rect 1078 171 1112 205
rect 1112 171 1150 205
rect 1150 171 1184 205
rect 1184 171 1222 205
rect 1222 171 1256 205
rect 1078 133 1256 171
rect 1078 99 1112 133
rect 1112 99 1150 133
rect 1150 99 1184 133
rect 1184 99 1222 133
rect 1222 99 1256 133
<< metal1 >>
rect 276 8166 1054 8172
rect 276 8132 288 8166
rect 322 8132 360 8166
rect 394 8132 432 8166
rect 466 8132 504 8166
rect 538 8132 576 8166
rect 610 8132 648 8166
rect 682 8132 720 8166
rect 754 8132 792 8166
rect 826 8132 864 8166
rect 898 8132 936 8166
rect 970 8132 1008 8166
rect 1042 8132 1054 8166
rect 276 8126 1054 8132
rect 68 8053 258 8065
rect 68 99 74 8053
rect 252 99 258 8053
rect 68 87 258 99
rect 1072 8053 1262 8065
rect 1072 99 1078 8053
rect 1256 99 1262 8053
rect 1072 87 1262 99
<< end >>
