magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< error_p >>
rect 111 372 117 378
rect 141 348 147 368
rect 183 260 189 280
rect 141 238 147 244
<< nwell >>
rect 0 309 352 630
<< pwell >>
rect 39 69 313 225
rect 69 31 103 69
<< scnmos >>
rect 117 95 147 199
rect 205 95 235 199
<< scpmoshvt >>
rect 117 387 147 545
rect 205 387 235 545
<< ndiff >>
rect 65 154 117 199
rect 65 120 73 154
rect 107 120 117 154
rect 65 95 117 120
rect 147 141 205 199
rect 147 107 159 141
rect 193 107 205 141
rect 147 95 205 107
rect 235 171 287 199
rect 235 137 245 171
rect 279 137 287 171
rect 235 95 287 137
<< pdiff >>
rect 65 525 117 545
rect 65 491 73 525
rect 107 491 117 525
rect 65 457 117 491
rect 65 423 73 457
rect 107 423 117 457
rect 65 387 117 423
rect 147 525 205 545
rect 147 491 159 525
rect 193 491 205 525
rect 147 457 205 491
rect 147 423 159 457
rect 193 423 205 457
rect 147 387 205 423
rect 235 525 287 545
rect 235 491 245 525
rect 279 491 287 525
rect 235 444 287 491
rect 235 410 245 444
rect 279 410 287 444
rect 235 387 287 410
<< ndiffc >>
rect 73 120 107 154
rect 159 107 193 141
rect 245 137 279 171
<< pdiffc >>
rect 73 491 107 525
rect 73 423 107 457
rect 159 491 193 525
rect 159 423 193 457
rect 245 491 279 525
rect 245 410 279 444
<< poly >>
rect 117 545 147 571
rect 205 545 235 571
rect 117 372 147 387
rect 111 348 147 372
rect 111 313 141 348
rect 205 326 235 387
rect 65 297 141 313
rect 65 263 75 297
rect 109 263 141 297
rect 65 247 141 263
rect 183 310 237 326
rect 183 276 193 310
rect 227 276 237 310
rect 183 260 237 276
rect 111 238 141 247
rect 111 214 147 238
rect 117 199 147 214
rect 205 199 235 260
rect 117 69 147 95
rect 205 69 235 95
<< polycont >>
rect 75 263 109 297
rect 193 276 227 310
<< locali >>
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 314 609
rect 71 525 107 541
rect 71 491 73 525
rect 71 457 107 491
rect 71 423 73 457
rect 143 525 209 575
rect 143 491 159 525
rect 193 491 209 525
rect 143 457 209 491
rect 143 423 159 457
rect 193 423 209 457
rect 243 525 297 541
rect 243 491 245 525
rect 279 491 297 525
rect 243 444 297 491
rect 71 389 107 423
rect 243 410 245 444
rect 279 410 297 444
rect 71 355 206 389
rect 243 360 297 410
rect 172 326 206 355
rect 59 297 127 319
rect 59 263 75 297
rect 109 263 127 297
rect 59 245 127 263
rect 172 310 227 326
rect 172 276 193 310
rect 172 260 227 276
rect 172 209 206 260
rect 73 175 206 209
rect 261 200 297 360
rect 73 154 107 175
rect 245 171 297 200
rect 73 99 107 120
rect 143 107 159 141
rect 193 107 209 141
rect 143 65 209 107
rect 279 137 297 171
rect 245 99 297 137
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 314 65
<< viali >>
rect 67 575 101 609
rect 159 575 193 609
rect 251 575 285 609
rect 67 31 101 65
rect 159 31 193 65
rect 251 31 285 65
<< metal1 >>
rect 38 609 314 640
rect 38 575 67 609
rect 101 575 159 609
rect 193 575 251 609
rect 285 575 314 609
rect 38 544 314 575
rect 38 65 314 96
rect 38 31 67 65
rect 101 31 159 65
rect 193 31 251 65
rect 285 31 314 65
rect 38 0 314 31
<< labels >>
flabel locali s 67 575 101 609 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
flabel locali s 69 31 103 65 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel locali s 249 133 283 167 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 249 405 283 439 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 249 473 283 507 0 FreeSans 200 0 0 0 X
port 6 nsew
flabel locali s 67 269 101 303 0 FreeSans 200 0 0 0 A
port 7 nsew
flabel pwell s 69 31 103 65 0 FreeSans 200 0 0 0 VNB
port 2 nsew
flabel nwell s 67 575 101 609 0 FreeSans 200 0 0 0 VPB
port 3 nsew
flabel metal1 s 69 31 103 65 0 FreeSans 200 0 0 0 VGND
port 4 nsew
flabel metal1 s 67 575 101 609 0 FreeSans 200 0 0 0 VPWR
port 5 nsew
rlabel comment s 38 48 38 48 4 buf_1
<< properties >>
string FIXED_BBOX 38 48 314 592
string path 0.190 2.960 1.570 2.960 
<< end >>
