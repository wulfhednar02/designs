magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -305 -380 7671 40720
<< l66d20 >>
rect 1020 -200 5020 40200
rect 1020 40200 5020 40530
<< l94d20 >>
rect -125 -125 6039 40125
<< l66d44 >>
rect 65 20275 235 20445
rect 425 20275 595 20445
rect 785 20275 955 20445
rect 5085 20275 5255 20445
rect 5445 20275 5615 20445
rect 5805 20275 5975 20445
rect 6258 20275 6428 20445
rect 6618 20275 6788 20445
rect 6978 20275 7148 20445
rect 65 30355 235 30525
rect 425 30355 595 30525
rect 785 30355 955 30525
rect 5085 30355 5255 30525
rect 5445 30355 5615 30525
rect 5805 30355 5975 30525
rect 6258 30355 6428 30525
rect 6618 30355 6788 30525
rect 6978 30355 7148 30525
rect 5085 35395 5255 35565
rect 5445 35395 5615 35565
rect 5805 35395 5975 35565
rect 6258 35395 6428 35565
rect 6618 35395 6788 35565
rect 6978 35395 7148 35565
rect 5445 37195 5615 37365
rect 5445 37555 5615 37725
rect 5445 37915 5615 38085
rect 5445 38275 5615 38445
rect 5445 38635 5615 38805
rect 5445 38995 5615 39165
rect 5445 39355 5615 39525
rect 5445 39715 5615 39885
rect 5445 35755 5615 35925
rect 5805 35755 5975 35925
rect 5805 36115 5975 36285
rect 5805 36475 5975 36645
rect 5805 36835 5975 37005
rect 5805 37195 5975 37365
rect 5805 37555 5975 37725
rect 5805 37915 5975 38085
rect 5805 38275 5975 38445
rect 5805 38635 5975 38805
rect 5805 38995 5975 39165
rect 5805 39355 5975 39525
rect 5805 39715 5975 39885
rect 5445 36115 5615 36285
rect 6258 35755 6428 35925
rect 6258 36115 6428 36285
rect 6258 36475 6428 36645
rect 6258 36835 6428 37005
rect 6258 37195 6428 37365
rect 6258 37555 6428 37725
rect 6258 37915 6428 38085
rect 6258 38275 6428 38445
rect 6258 38635 6428 38805
rect 6258 38995 6428 39165
rect 6258 39355 6428 39525
rect 6258 39715 6428 39885
rect 5445 36475 5615 36645
rect 6618 35755 6788 35925
rect 6618 36115 6788 36285
rect 6618 36475 6788 36645
rect 6618 36835 6788 37005
rect 6618 37195 6788 37365
rect 6618 37555 6788 37725
rect 6618 37915 6788 38085
rect 6618 38275 6788 38445
rect 6618 38635 6788 38805
rect 6618 38995 6788 39165
rect 6618 39355 6788 39525
rect 6618 39715 6788 39885
rect 5445 36835 5615 37005
rect 6978 35755 7148 35925
rect 6978 36115 7148 36285
rect 6978 36475 7148 36645
rect 6978 36835 7148 37005
rect 6978 37195 7148 37365
rect 6978 37555 7148 37725
rect 6978 37915 7148 38085
rect 6978 38275 7148 38445
rect 6978 38635 7148 38805
rect 6978 38995 7148 39165
rect 6978 39355 7148 39525
rect 6978 39715 7148 39885
rect 5085 38995 5255 39165
rect 5085 39355 5255 39525
rect 5085 39715 5255 39885
rect 5085 35755 5255 35925
rect 5085 36115 5255 36285
rect 3655 40280 3825 40450
rect 4015 40280 4185 40450
rect 4375 40280 4545 40450
rect 4735 40280 4905 40450
rect 5085 36475 5255 36645
rect 5085 36835 5255 37005
rect 5085 37195 5255 37365
rect 5085 37555 5255 37725
rect 5085 37915 5255 38085
rect 5085 38275 5255 38445
rect 5085 38635 5255 38805
rect 5085 32875 5255 33045
rect 5085 33235 5255 33405
rect 5085 33595 5255 33765
rect 5085 33955 5255 34125
rect 5085 30715 5255 30885
rect 5085 34315 5255 34485
rect 5085 34675 5255 34845
rect 5085 31435 5255 31605
rect 5085 35035 5255 35205
rect 5085 32515 5255 32685
rect 5085 31795 5255 31965
rect 5085 31075 5255 31245
rect 5085 32155 5255 32325
rect 5805 33235 5975 33405
rect 5805 33595 5975 33765
rect 5805 33955 5975 34125
rect 5805 34315 5975 34485
rect 5805 34675 5975 34845
rect 5805 35035 5975 35205
rect 5445 31075 5615 31245
rect 5445 31435 5615 31605
rect 5445 31795 5615 31965
rect 5445 32155 5615 32325
rect 5445 32515 5615 32685
rect 5445 32875 5615 33045
rect 6618 30715 6788 30885
rect 6618 31075 6788 31245
rect 6618 31435 6788 31605
rect 6618 31795 6788 31965
rect 6618 32155 6788 32325
rect 6618 32515 6788 32685
rect 6618 32875 6788 33045
rect 6618 33235 6788 33405
rect 6618 33595 6788 33765
rect 6618 33955 6788 34125
rect 6618 34315 6788 34485
rect 6618 34675 6788 34845
rect 6618 35035 6788 35205
rect 5445 33235 5615 33405
rect 5445 33595 5615 33765
rect 5445 33955 5615 34125
rect 5445 34315 5615 34485
rect 5445 34675 5615 34845
rect 5445 35035 5615 35205
rect 5445 30715 5615 30885
rect 5805 30715 5975 30885
rect 5805 31075 5975 31245
rect 5805 31435 5975 31605
rect 5805 31795 5975 31965
rect 5805 32155 5975 32325
rect 6258 30715 6428 30885
rect 6258 31075 6428 31245
rect 6978 30715 7148 30885
rect 6978 31075 7148 31245
rect 6978 31435 7148 31605
rect 6978 31795 7148 31965
rect 6978 32155 7148 32325
rect 6978 32515 7148 32685
rect 6978 32875 7148 33045
rect 6978 33235 7148 33405
rect 6978 33595 7148 33765
rect 6978 33955 7148 34125
rect 6978 34315 7148 34485
rect 6978 34675 7148 34845
rect 6978 35035 7148 35205
rect 6258 31435 6428 31605
rect 6258 31795 6428 31965
rect 6258 32155 6428 32325
rect 6258 32515 6428 32685
rect 6258 32875 6428 33045
rect 6258 33235 6428 33405
rect 6258 33595 6428 33765
rect 6258 33955 6428 34125
rect 6258 34315 6428 34485
rect 6258 34675 6428 34845
rect 6258 35035 6428 35205
rect 5805 32515 5975 32685
rect 5805 32875 5975 33045
rect 65 32515 235 32685
rect 65 32875 235 33045
rect 65 33235 235 33405
rect 65 33595 235 33765
rect 65 33955 235 34125
rect 65 34315 235 34485
rect 65 34675 235 34845
rect 65 35035 235 35205
rect 65 35395 235 35565
rect 65 35755 235 35925
rect 65 36115 235 36285
rect 65 36475 235 36645
rect 65 36835 235 37005
rect 65 37195 235 37365
rect 65 37555 235 37725
rect 65 37915 235 38085
rect 65 38275 235 38445
rect 65 38635 235 38805
rect 65 38995 235 39165
rect 65 39355 235 39525
rect 65 39715 235 39885
rect 65 30715 235 30885
rect 425 30715 595 30885
rect 425 31075 595 31245
rect 425 31435 595 31605
rect 425 31795 595 31965
rect 425 32155 595 32325
rect 425 32515 595 32685
rect 425 32875 595 33045
rect 425 33235 595 33405
rect 425 33595 595 33765
rect 425 33955 595 34125
rect 425 34315 595 34485
rect 425 34675 595 34845
rect 425 35035 595 35205
rect 425 35395 595 35565
rect 425 35755 595 35925
rect 425 36115 595 36285
rect 425 36475 595 36645
rect 425 36835 595 37005
rect 425 37195 595 37365
rect 425 37555 595 37725
rect 425 37915 595 38085
rect 425 38275 595 38445
rect 425 38635 595 38805
rect 425 38995 595 39165
rect 425 39355 595 39525
rect 425 39715 595 39885
rect 65 31075 235 31245
rect 785 30715 955 30885
rect 785 31075 955 31245
rect 785 31435 955 31605
rect 785 31795 955 31965
rect 785 32155 955 32325
rect 785 32515 955 32685
rect 785 32875 955 33045
rect 785 33235 955 33405
rect 785 33595 955 33765
rect 785 33955 955 34125
rect 785 34315 955 34485
rect 785 34675 955 34845
rect 785 35035 955 35205
rect 785 35395 955 35565
rect 785 35755 955 35925
rect 785 36115 955 36285
rect 785 36475 955 36645
rect 785 36835 955 37005
rect 785 37195 955 37365
rect 785 37555 955 37725
rect 785 37915 955 38085
rect 785 38275 955 38445
rect 785 38635 955 38805
rect 785 38995 955 39165
rect 785 39355 955 39525
rect 785 39715 955 39885
rect 65 31435 235 31605
rect 65 31795 235 31965
rect 65 32155 235 32325
rect 1135 40280 1305 40450
rect 1495 40280 1665 40450
rect 1855 40280 2025 40450
rect 2215 40280 2385 40450
rect 2575 40280 2745 40450
rect 2935 40280 3105 40450
rect 3295 40280 3465 40450
rect 425 22435 595 22605
rect 425 22795 595 22965
rect 65 20995 235 21165
rect 785 20635 955 20805
rect 785 20995 955 21165
rect 785 21355 955 21525
rect 785 21715 955 21885
rect 785 22075 955 22245
rect 785 22435 955 22605
rect 65 21715 235 21885
rect 785 22795 955 22965
rect 785 23155 955 23325
rect 785 23515 955 23685
rect 785 23875 955 24045
rect 785 24235 955 24405
rect 785 24595 955 24765
rect 785 24955 955 25125
rect 785 25315 955 25485
rect 785 25675 955 25845
rect 785 26035 955 26205
rect 785 26395 955 26565
rect 785 26755 955 26925
rect 785 27115 955 27285
rect 785 27475 955 27645
rect 785 27835 955 28005
rect 65 22795 235 22965
rect 785 28195 955 28365
rect 785 28555 955 28725
rect 785 28915 955 29085
rect 785 29275 955 29445
rect 785 29635 955 29805
rect 785 29995 955 30165
rect 425 23155 595 23325
rect 425 23515 595 23685
rect 425 23875 595 24045
rect 425 24235 595 24405
rect 425 24595 595 24765
rect 425 24955 595 25125
rect 65 22075 235 22245
rect 425 25315 595 25485
rect 425 25675 595 25845
rect 425 26035 595 26205
rect 425 26395 595 26565
rect 425 26755 595 26925
rect 425 27115 595 27285
rect 425 27475 595 27645
rect 425 27835 595 28005
rect 425 28195 595 28365
rect 425 28555 595 28725
rect 425 28915 595 29085
rect 425 29275 595 29445
rect 425 29635 595 29805
rect 425 29995 595 30165
rect 65 23155 235 23325
rect 65 26395 235 26565
rect 65 26755 235 26925
rect 65 27115 235 27285
rect 65 27475 235 27645
rect 65 27835 235 28005
rect 65 28195 235 28365
rect 65 28555 235 28725
rect 65 21355 235 21525
rect 65 28915 235 29085
rect 65 29275 235 29445
rect 65 29635 235 29805
rect 65 29995 235 30165
rect 65 23515 235 23685
rect 65 23875 235 24045
rect 65 24235 235 24405
rect 65 24595 235 24765
rect 65 24955 235 25125
rect 65 25315 235 25485
rect 65 25675 235 25845
rect 65 26035 235 26205
rect 65 20635 235 20805
rect 425 20635 595 20805
rect 425 20995 595 21165
rect 425 21355 595 21525
rect 65 22435 235 22605
rect 425 21715 595 21885
rect 425 22075 595 22245
rect 6258 25315 6428 25485
rect 6618 25315 6788 25485
rect 5805 25315 5975 25485
rect 5445 25315 5615 25485
rect 6978 25315 7148 25485
rect 5085 25315 5255 25485
rect 6258 27475 6428 27645
rect 6258 27835 6428 28005
rect 6258 28195 6428 28365
rect 6258 28555 6428 28725
rect 6258 28915 6428 29085
rect 6258 29275 6428 29445
rect 6258 29635 6428 29805
rect 6258 29995 6428 30165
rect 6258 25675 6428 25845
rect 6618 25675 6788 25845
rect 6618 26035 6788 26205
rect 6618 26395 6788 26565
rect 6618 26755 6788 26925
rect 6618 27115 6788 27285
rect 6618 27475 6788 27645
rect 6618 27835 6788 28005
rect 6618 28195 6788 28365
rect 6618 28555 6788 28725
rect 6618 28915 6788 29085
rect 6618 29275 6788 29445
rect 6618 29635 6788 29805
rect 6618 29995 6788 30165
rect 6258 26035 6428 26205
rect 5805 25675 5975 25845
rect 5805 26035 5975 26205
rect 5805 26395 5975 26565
rect 5805 26755 5975 26925
rect 5805 27115 5975 27285
rect 5805 27475 5975 27645
rect 5805 27835 5975 28005
rect 5805 28195 5975 28365
rect 5805 28555 5975 28725
rect 5805 28915 5975 29085
rect 5805 29275 5975 29445
rect 5805 29635 5975 29805
rect 5805 29995 5975 30165
rect 6258 26395 6428 26565
rect 5445 25675 5615 25845
rect 6258 26755 6428 26925
rect 6978 25675 7148 25845
rect 6978 26035 7148 26205
rect 6978 26395 7148 26565
rect 6978 26755 7148 26925
rect 6978 27115 7148 27285
rect 6978 27475 7148 27645
rect 6978 27835 7148 28005
rect 6978 28195 7148 28365
rect 6978 28555 7148 28725
rect 6978 28915 7148 29085
rect 6978 29275 7148 29445
rect 6978 29635 7148 29805
rect 6978 29995 7148 30165
rect 5445 26035 5615 26205
rect 5445 26395 5615 26565
rect 5445 26755 5615 26925
rect 5445 27115 5615 27285
rect 5445 27475 5615 27645
rect 5445 27835 5615 28005
rect 5445 28195 5615 28365
rect 5445 28555 5615 28725
rect 5445 28915 5615 29085
rect 5445 29275 5615 29445
rect 5445 29635 5615 29805
rect 5445 29995 5615 30165
rect 6258 27115 6428 27285
rect 5085 27475 5255 27645
rect 5085 27835 5255 28005
rect 5085 28195 5255 28365
rect 5085 28555 5255 28725
rect 5085 28915 5255 29085
rect 5085 29275 5255 29445
rect 5085 29635 5255 29805
rect 5085 29995 5255 30165
rect 5085 25675 5255 25845
rect 5085 26035 5255 26205
rect 5085 26395 5255 26565
rect 5085 26755 5255 26925
rect 5085 27115 5255 27285
rect 5085 20995 5255 21165
rect 5085 21355 5255 21525
rect 5085 21715 5255 21885
rect 5085 22075 5255 22245
rect 5085 22435 5255 22605
rect 5085 22795 5255 22965
rect 5085 23155 5255 23325
rect 5085 23515 5255 23685
rect 5085 23875 5255 24045
rect 5085 24235 5255 24405
rect 5085 24595 5255 24765
rect 5085 24955 5255 25125
rect 5085 20635 5255 20805
rect 5445 22075 5615 22245
rect 5445 22435 5615 22605
rect 5445 22795 5615 22965
rect 5445 23155 5615 23325
rect 5445 23515 5615 23685
rect 5445 23875 5615 24045
rect 5445 24235 5615 24405
rect 5445 24595 5615 24765
rect 5445 24955 5615 25125
rect 6618 21715 6788 21885
rect 6618 22075 6788 22245
rect 6978 20635 7148 20805
rect 6978 20995 7148 21165
rect 6978 21355 7148 21525
rect 6978 21715 7148 21885
rect 6978 22075 7148 22245
rect 6978 22435 7148 22605
rect 6978 22795 7148 22965
rect 6978 23155 7148 23325
rect 6978 23515 7148 23685
rect 6978 23875 7148 24045
rect 6978 24235 7148 24405
rect 6978 24595 7148 24765
rect 6978 24955 7148 25125
rect 6618 22435 6788 22605
rect 6618 22795 6788 22965
rect 6618 23155 6788 23325
rect 6618 23515 6788 23685
rect 6618 23875 6788 24045
rect 6618 24235 6788 24405
rect 6618 24595 6788 24765
rect 6618 24955 6788 25125
rect 6258 23515 6428 23685
rect 6258 23875 6428 24045
rect 6258 24235 6428 24405
rect 6258 24595 6428 24765
rect 6258 24955 6428 25125
rect 6258 21355 6428 21525
rect 6258 21715 6428 21885
rect 6258 22075 6428 22245
rect 6258 22435 6428 22605
rect 6258 22795 6428 22965
rect 6258 23155 6428 23325
rect 5445 20635 5615 20805
rect 5805 20635 5975 20805
rect 5805 20995 5975 21165
rect 5805 21355 5975 21525
rect 5805 21715 5975 21885
rect 5805 22075 5975 22245
rect 5805 22435 5975 22605
rect 5805 22795 5975 22965
rect 5805 23155 5975 23325
rect 5805 23515 5975 23685
rect 5805 23875 5975 24045
rect 5805 24235 5975 24405
rect 5805 24595 5975 24765
rect 5805 24955 5975 25125
rect 6618 20635 6788 20805
rect 6618 20995 6788 21165
rect 6618 21355 6788 21525
rect 5445 20995 5615 21165
rect 5445 21355 5615 21525
rect 5445 21715 5615 21885
rect 6258 20635 6428 20805
rect 6258 20995 6428 21165
rect 785 10195 955 10365
rect 5805 10195 5975 10365
rect 425 10195 595 10365
rect 6258 10195 6428 10365
rect 5085 10195 5255 10365
rect 6618 10195 6788 10365
rect 65 10195 235 10365
rect 6978 10195 7148 10365
rect 5445 10195 5615 10365
rect 5805 15235 5975 15405
rect 6258 15235 6428 15405
rect 5085 15235 5255 15405
rect 6618 15235 6788 15405
rect 6978 15235 7148 15405
rect 5445 15235 5615 15405
rect 5805 17395 5975 17565
rect 5805 17755 5975 17925
rect 5805 18115 5975 18285
rect 5805 18475 5975 18645
rect 5805 18835 5975 19005
rect 5805 19195 5975 19365
rect 5805 19555 5975 19725
rect 5805 19915 5975 20085
rect 5805 15595 5975 15765
rect 6258 15595 6428 15765
rect 6258 15955 6428 16125
rect 6258 16315 6428 16485
rect 6258 16675 6428 16845
rect 6258 17035 6428 17205
rect 6258 17395 6428 17565
rect 6258 17755 6428 17925
rect 6258 18115 6428 18285
rect 6258 18475 6428 18645
rect 6258 18835 6428 19005
rect 6258 19195 6428 19365
rect 6258 19555 6428 19725
rect 6258 19915 6428 20085
rect 5805 15955 5975 16125
rect 5805 16315 5975 16485
rect 6618 15595 6788 15765
rect 6618 15955 6788 16125
rect 6618 16315 6788 16485
rect 6618 16675 6788 16845
rect 6618 17035 6788 17205
rect 6618 17395 6788 17565
rect 6618 17755 6788 17925
rect 6618 18115 6788 18285
rect 6618 18475 6788 18645
rect 6618 18835 6788 19005
rect 6618 19195 6788 19365
rect 6618 19555 6788 19725
rect 6618 19915 6788 20085
rect 5805 16675 5975 16845
rect 6978 15595 7148 15765
rect 6978 15955 7148 16125
rect 6978 16315 7148 16485
rect 6978 16675 7148 16845
rect 6978 17035 7148 17205
rect 6978 17395 7148 17565
rect 6978 17755 7148 17925
rect 6978 18115 7148 18285
rect 6978 18475 7148 18645
rect 6978 18835 7148 19005
rect 6978 19195 7148 19365
rect 6978 19555 7148 19725
rect 6978 19915 7148 20085
rect 5805 17035 5975 17205
rect 5445 15595 5615 15765
rect 5445 15955 5615 16125
rect 5445 16315 5615 16485
rect 5445 16675 5615 16845
rect 5445 17035 5615 17205
rect 5445 17395 5615 17565
rect 5445 17755 5615 17925
rect 5445 18115 5615 18285
rect 5445 18475 5615 18645
rect 5445 18835 5615 19005
rect 5445 19195 5615 19365
rect 5445 19555 5615 19725
rect 5445 19915 5615 20085
rect 5085 16675 5255 16845
rect 5085 17035 5255 17205
rect 5085 17395 5255 17565
rect 5085 17755 5255 17925
rect 5085 18115 5255 18285
rect 5085 18475 5255 18645
rect 5085 18835 5255 19005
rect 5085 19195 5255 19365
rect 5085 19555 5255 19725
rect 5085 19915 5255 20085
rect 5085 15595 5255 15765
rect 5085 15955 5255 16125
rect 5085 16315 5255 16485
rect 5085 11995 5255 12165
rect 5085 12355 5255 12525
rect 5085 12715 5255 12885
rect 5085 13075 5255 13245
rect 5085 13435 5255 13605
rect 5085 13795 5255 13965
rect 5085 14155 5255 14325
rect 5085 14515 5255 14685
rect 5085 14875 5255 15045
rect 5085 10555 5255 10725
rect 5085 10915 5255 11085
rect 5085 11275 5255 11445
rect 5085 11635 5255 11805
rect 5805 13075 5975 13245
rect 5805 13435 5975 13605
rect 5805 10555 5975 10725
rect 5805 10915 5975 11085
rect 6258 10555 6428 10725
rect 6258 10915 6428 11085
rect 6258 11275 6428 11445
rect 6258 11635 6428 11805
rect 5805 11995 5975 12165
rect 5805 12355 5975 12525
rect 6978 10555 7148 10725
rect 6978 10915 7148 11085
rect 6978 11275 7148 11445
rect 6978 11635 7148 11805
rect 6978 11995 7148 12165
rect 6978 12355 7148 12525
rect 6978 12715 7148 12885
rect 6978 13075 7148 13245
rect 6978 13435 7148 13605
rect 6978 13795 7148 13965
rect 6978 14155 7148 14325
rect 6978 14515 7148 14685
rect 6978 14875 7148 15045
rect 6258 11995 6428 12165
rect 6258 12355 6428 12525
rect 5805 11275 5975 11445
rect 6258 12715 6428 12885
rect 6258 13075 6428 13245
rect 6258 13435 6428 13605
rect 6258 13795 6428 13965
rect 6258 14155 6428 14325
rect 5805 11635 5975 11805
rect 6618 10555 6788 10725
rect 6618 10915 6788 11085
rect 6618 11275 6788 11445
rect 6618 11635 6788 11805
rect 6618 11995 6788 12165
rect 5805 12715 5975 12885
rect 5445 10555 5615 10725
rect 5445 10915 5615 11085
rect 5445 11275 5615 11445
rect 5445 11635 5615 11805
rect 5445 11995 5615 12165
rect 5445 12355 5615 12525
rect 5445 12715 5615 12885
rect 5445 13075 5615 13245
rect 5445 13435 5615 13605
rect 5445 13795 5615 13965
rect 5445 14155 5615 14325
rect 5445 14515 5615 14685
rect 5445 14875 5615 15045
rect 6618 12355 6788 12525
rect 6618 12715 6788 12885
rect 6618 13075 6788 13245
rect 6618 13435 6788 13605
rect 6618 13795 6788 13965
rect 6618 14155 6788 14325
rect 6618 14515 6788 14685
rect 6618 14875 6788 15045
rect 6258 14515 6428 14685
rect 6258 14875 6428 15045
rect 5805 13795 5975 13965
rect 5805 14155 5975 14325
rect 5805 14515 5975 14685
rect 5805 14875 5975 15045
rect 65 10555 235 10725
rect 65 10915 235 11085
rect 65 11275 235 11445
rect 65 11635 235 11805
rect 65 11995 235 12165
rect 65 12355 235 12525
rect 65 12715 235 12885
rect 65 13075 235 13245
rect 65 13435 235 13605
rect 65 13795 235 13965
rect 65 14155 235 14325
rect 65 14515 235 14685
rect 65 14875 235 15045
rect 65 15235 235 15405
rect 65 15595 235 15765
rect 65 15955 235 16125
rect 65 16315 235 16485
rect 65 16675 235 16845
rect 65 17035 235 17205
rect 65 17395 235 17565
rect 65 17755 235 17925
rect 65 18115 235 18285
rect 65 18475 235 18645
rect 425 11995 595 12165
rect 425 12355 595 12525
rect 425 12715 595 12885
rect 425 13075 595 13245
rect 425 13435 595 13605
rect 425 13795 595 13965
rect 425 14155 595 14325
rect 425 14515 595 14685
rect 425 14875 595 15045
rect 425 15235 595 15405
rect 425 15595 595 15765
rect 425 15955 595 16125
rect 425 16315 595 16485
rect 425 16675 595 16845
rect 425 17035 595 17205
rect 425 17395 595 17565
rect 425 17755 595 17925
rect 425 18115 595 18285
rect 425 18475 595 18645
rect 425 18835 595 19005
rect 425 19195 595 19365
rect 785 12355 955 12525
rect 785 12715 955 12885
rect 785 13075 955 13245
rect 425 19555 595 19725
rect 425 19915 595 20085
rect 65 19915 235 20085
rect 785 13435 955 13605
rect 785 13795 955 13965
rect 785 14155 955 14325
rect 785 14515 955 14685
rect 785 14875 955 15045
rect 785 15235 955 15405
rect 785 15595 955 15765
rect 785 15955 955 16125
rect 785 16315 955 16485
rect 785 16675 955 16845
rect 785 17035 955 17205
rect 785 17395 955 17565
rect 785 17755 955 17925
rect 785 18115 955 18285
rect 785 18475 955 18645
rect 785 18835 955 19005
rect 785 10555 955 10725
rect 785 10915 955 11085
rect 785 11275 955 11445
rect 785 11635 955 11805
rect 785 19195 955 19365
rect 785 19555 955 19725
rect 785 19915 955 20085
rect 65 19555 235 19725
rect 785 11995 955 12165
rect 425 10555 595 10725
rect 425 10915 595 11085
rect 425 11275 595 11445
rect 425 11635 595 11805
rect 65 18835 235 19005
rect 65 19195 235 19365
rect 785 8755 955 8925
rect 785 9115 955 9285
rect 785 9475 955 9645
rect 785 9835 955 10005
rect 785 1555 955 1725
rect 785 1915 955 2085
rect 785 2275 955 2445
rect 785 2635 955 2805
rect 785 2995 955 3165
rect 785 3355 955 3525
rect 785 3715 955 3885
rect 785 4075 955 4245
rect 785 4435 955 4605
rect 425 115 595 285
rect 425 475 595 645
rect 425 835 595 1005
rect 425 1195 595 1365
rect 425 1555 595 1725
rect 425 1915 595 2085
rect 425 2275 595 2445
rect 425 2635 595 2805
rect 425 2995 595 3165
rect 65 115 235 285
rect 65 475 235 645
rect 65 835 235 1005
rect 65 1195 235 1365
rect 425 3355 595 3525
rect 425 3715 595 3885
rect 425 4075 595 4245
rect 425 4435 595 4605
rect 425 4795 595 4965
rect 425 5155 595 5325
rect 425 5515 595 5685
rect 425 5875 595 6045
rect 425 6235 595 6405
rect 425 6595 595 6765
rect 425 6955 595 7125
rect 425 7315 595 7485
rect 425 7675 595 7845
rect 425 8035 595 8205
rect 425 8395 595 8565
rect 425 8755 595 8925
rect 425 9115 595 9285
rect 425 9475 595 9645
rect 425 9835 595 10005
rect 785 4795 955 4965
rect 785 5155 955 5325
rect 785 5515 955 5685
rect 785 5875 955 6045
rect 785 6235 955 6405
rect 785 6595 955 6765
rect 785 6955 955 7125
rect 785 7315 955 7485
rect 785 7675 955 7845
rect 65 1555 235 1725
rect 65 1915 235 2085
rect 65 2275 235 2445
rect 65 2635 235 2805
rect 65 2995 235 3165
rect 65 3355 235 3525
rect 65 3715 235 3885
rect 65 4075 235 4245
rect 65 4435 235 4605
rect 65 4795 235 4965
rect 65 5155 235 5325
rect 65 5515 235 5685
rect 65 5875 235 6045
rect 65 6235 235 6405
rect 65 6595 235 6765
rect 65 6955 235 7125
rect 65 7315 235 7485
rect 65 7675 235 7845
rect 65 8035 235 8205
rect 65 8395 235 8565
rect 65 8755 235 8925
rect 65 9115 235 9285
rect 65 9475 235 9645
rect 65 9835 235 10005
rect 785 8035 955 8205
rect 785 8395 955 8565
rect 785 115 955 285
rect 785 475 955 645
rect 785 835 955 1005
rect 785 1195 955 1365
rect 5085 5155 5255 5325
rect 6258 5155 6428 5325
rect 6978 5155 7148 5325
rect 6618 5155 6788 5325
rect 5445 5155 5615 5325
rect 5805 5155 5975 5325
rect 6258 6595 6428 6765
rect 5805 9835 5975 10005
rect 6978 5515 7148 5685
rect 6978 5875 7148 6045
rect 6978 6235 7148 6405
rect 6978 6595 7148 6765
rect 6978 6955 7148 7125
rect 6978 7315 7148 7485
rect 6978 7675 7148 7845
rect 6978 8035 7148 8205
rect 6978 8395 7148 8565
rect 6978 8755 7148 8925
rect 6978 9115 7148 9285
rect 6978 9475 7148 9645
rect 6978 9835 7148 10005
rect 6258 6955 6428 7125
rect 6258 7315 6428 7485
rect 6258 7675 6428 7845
rect 6258 8035 6428 8205
rect 6258 8395 6428 8565
rect 6258 8755 6428 8925
rect 6258 9115 6428 9285
rect 6258 9475 6428 9645
rect 6258 5515 6428 5685
rect 6618 5515 6788 5685
rect 6618 5875 6788 6045
rect 6618 6235 6788 6405
rect 6618 6595 6788 6765
rect 6618 6955 6788 7125
rect 6258 5875 6428 6045
rect 5445 5515 5615 5685
rect 5445 5875 5615 6045
rect 5445 6235 5615 6405
rect 5445 6595 5615 6765
rect 5445 6955 5615 7125
rect 5445 7315 5615 7485
rect 5445 7675 5615 7845
rect 5445 8035 5615 8205
rect 5445 8395 5615 8565
rect 5445 8755 5615 8925
rect 5445 9115 5615 9285
rect 5445 9475 5615 9645
rect 5445 9835 5615 10005
rect 6618 7315 6788 7485
rect 6618 7675 6788 7845
rect 6618 8035 6788 8205
rect 6618 8395 6788 8565
rect 6618 8755 6788 8925
rect 6618 9115 6788 9285
rect 6618 9475 6788 9645
rect 6618 9835 6788 10005
rect 6258 9835 6428 10005
rect 6258 6235 6428 6405
rect 5805 5515 5975 5685
rect 5805 5875 5975 6045
rect 5805 6235 5975 6405
rect 5805 6595 5975 6765
rect 5805 6955 5975 7125
rect 5805 7315 5975 7485
rect 5805 7675 5975 7845
rect 5805 8035 5975 8205
rect 5805 8395 5975 8565
rect 5805 8755 5975 8925
rect 5805 9115 5975 9285
rect 5805 9475 5975 9645
rect 5085 6955 5255 7125
rect 5085 7315 5255 7485
rect 5085 7675 5255 7845
rect 5085 8035 5255 8205
rect 5085 8395 5255 8565
rect 5085 8755 5255 8925
rect 5085 9115 5255 9285
rect 5085 9475 5255 9645
rect 5085 9835 5255 10005
rect 5085 5515 5255 5685
rect 5085 5875 5255 6045
rect 5085 6235 5255 6405
rect 5085 6595 5255 6765
rect 5085 2635 5255 2805
rect 5085 3715 5255 3885
rect 5085 4075 5255 4245
rect 5085 4435 5255 4605
rect 5085 4795 5255 4965
rect 5085 2995 5255 3165
rect 5085 3355 5255 3525
rect 5085 115 5255 285
rect 5085 475 5255 645
rect 5085 835 5255 1005
rect 5085 1195 5255 1365
rect 5085 1555 5255 1725
rect 5085 1915 5255 2085
rect 5085 2275 5255 2445
rect 6618 1915 6788 2085
rect 6618 2275 6788 2445
rect 6618 2635 6788 2805
rect 6618 2995 6788 3165
rect 6618 3355 6788 3525
rect 6618 3715 6788 3885
rect 6618 4075 6788 4245
rect 6618 4435 6788 4605
rect 6618 4795 6788 4965
rect 5445 2275 5615 2445
rect 6978 115 7148 285
rect 6978 475 7148 645
rect 6978 835 7148 1005
rect 6978 1195 7148 1365
rect 6978 1555 7148 1725
rect 5445 2635 5615 2805
rect 5445 2995 5615 3165
rect 5445 3355 5615 3525
rect 5445 3715 5615 3885
rect 5445 4075 5615 4245
rect 5445 4435 5615 4605
rect 5445 4795 5615 4965
rect 6978 1915 7148 2085
rect 6978 2275 7148 2445
rect 6978 2635 7148 2805
rect 6978 2995 7148 3165
rect 6978 3355 7148 3525
rect 6978 3715 7148 3885
rect 6978 4075 7148 4245
rect 6978 4435 7148 4605
rect 6978 4795 7148 4965
rect 6258 1195 6428 1365
rect 6258 1555 6428 1725
rect 6258 1915 6428 2085
rect 6258 2275 6428 2445
rect 6258 2635 6428 2805
rect 6258 2995 6428 3165
rect 6258 3355 6428 3525
rect 6258 3715 6428 3885
rect 6258 4075 6428 4245
rect 6258 4435 6428 4605
rect 6258 4795 6428 4965
rect 5805 115 5975 285
rect 5805 475 5975 645
rect 6258 115 6428 285
rect 5805 835 5975 1005
rect 5805 1195 5975 1365
rect 5805 1555 5975 1725
rect 5805 1915 5975 2085
rect 5805 2275 5975 2445
rect 5805 2635 5975 2805
rect 5805 2995 5975 3165
rect 5805 3355 5975 3525
rect 5805 3715 5975 3885
rect 5805 4075 5975 4245
rect 5805 4435 5975 4605
rect 5805 4795 5975 4965
rect 6258 475 6428 645
rect 6258 835 6428 1005
rect 5445 115 5615 285
rect 5445 475 5615 645
rect 5445 835 5615 1005
rect 5445 1195 5615 1365
rect 5445 1555 5615 1725
rect 5445 1915 5615 2085
rect 6618 115 6788 285
rect 6618 475 6788 645
rect 6618 835 6788 1005
rect 6618 1195 6788 1365
rect 6618 1555 6788 1725
<< l67d44 >>
rect 65 20275 235 20445
rect 425 20275 595 20445
rect 785 20275 955 20445
rect 5085 20275 5255 20445
rect 5445 20275 5615 20445
rect 5805 20275 5975 20445
rect 65 30355 235 30525
rect 425 30355 595 30525
rect 785 30355 955 30525
rect 5085 30355 5255 30525
rect 5445 30355 5615 30525
rect 5805 30355 5975 30525
rect 2935 40280 3105 40450
rect 5085 31795 5255 31965
rect 5085 32155 5255 32325
rect 5085 32515 5255 32685
rect 5085 32875 5255 33045
rect 5085 33235 5255 33405
rect 5085 33595 5255 33765
rect 5085 33955 5255 34125
rect 5085 34315 5255 34485
rect 5085 34675 5255 34845
rect 5085 35035 5255 35205
rect 5085 35395 5255 35565
rect 5085 35755 5255 35925
rect 5085 36115 5255 36285
rect 5085 36475 5255 36645
rect 5085 36835 5255 37005
rect 5085 37195 5255 37365
rect 5085 37555 5255 37725
rect 5085 37915 5255 38085
rect 5085 38275 5255 38445
rect 5085 38635 5255 38805
rect 5085 38995 5255 39165
rect 5085 39355 5255 39525
rect 5085 39715 5255 39885
rect 5085 30715 5255 30885
rect 5445 30715 5615 30885
rect 5445 31075 5615 31245
rect 5445 31435 5615 31605
rect 5445 31795 5615 31965
rect 5445 32155 5615 32325
rect 5445 32515 5615 32685
rect 5445 32875 5615 33045
rect 5445 33235 5615 33405
rect 5445 33595 5615 33765
rect 5445 33955 5615 34125
rect 5445 34315 5615 34485
rect 5445 34675 5615 34845
rect 5445 35035 5615 35205
rect 5445 35395 5615 35565
rect 5445 35755 5615 35925
rect 5445 36115 5615 36285
rect 5445 36475 5615 36645
rect 5445 36835 5615 37005
rect 5445 37195 5615 37365
rect 5445 37555 5615 37725
rect 5445 37915 5615 38085
rect 5445 38275 5615 38445
rect 5445 38635 5615 38805
rect 5445 38995 5615 39165
rect 5445 39355 5615 39525
rect 5445 39715 5615 39885
rect 5085 31075 5255 31245
rect 5805 30715 5975 30885
rect 5805 31075 5975 31245
rect 5805 31435 5975 31605
rect 5805 31795 5975 31965
rect 5805 32155 5975 32325
rect 5805 32515 5975 32685
rect 5805 32875 5975 33045
rect 5805 33235 5975 33405
rect 5805 33595 5975 33765
rect 5805 33955 5975 34125
rect 5805 34315 5975 34485
rect 5805 34675 5975 34845
rect 5805 35035 5975 35205
rect 5805 35395 5975 35565
rect 5805 35755 5975 35925
rect 5805 36115 5975 36285
rect 5805 36475 5975 36645
rect 5805 36835 5975 37005
rect 5805 37195 5975 37365
rect 5805 37555 5975 37725
rect 5805 37915 5975 38085
rect 5805 38275 5975 38445
rect 5805 38635 5975 38805
rect 5805 38995 5975 39165
rect 5805 39355 5975 39525
rect 5805 39715 5975 39885
rect 5085 31435 5255 31605
rect 3295 40280 3465 40450
rect 3655 40280 3825 40450
rect 4015 40280 4185 40450
rect 4375 40280 4545 40450
rect 4735 40280 4905 40450
rect 65 34675 235 34845
rect 65 35035 235 35205
rect 65 35395 235 35565
rect 65 35755 235 35925
rect 65 36115 235 36285
rect 65 36475 235 36645
rect 65 36835 235 37005
rect 65 37195 235 37365
rect 65 37555 235 37725
rect 65 37915 235 38085
rect 65 38275 235 38445
rect 65 38635 235 38805
rect 65 38995 235 39165
rect 65 39355 235 39525
rect 65 39715 235 39885
rect 65 30715 235 30885
rect 425 30715 595 30885
rect 425 31075 595 31245
rect 425 31435 595 31605
rect 425 31795 595 31965
rect 425 32155 595 32325
rect 425 32515 595 32685
rect 425 32875 595 33045
rect 425 33235 595 33405
rect 425 33595 595 33765
rect 425 33955 595 34125
rect 425 34315 595 34485
rect 425 34675 595 34845
rect 425 35035 595 35205
rect 425 35395 595 35565
rect 425 35755 595 35925
rect 425 36115 595 36285
rect 425 36475 595 36645
rect 425 36835 595 37005
rect 425 37195 595 37365
rect 425 37555 595 37725
rect 425 37915 595 38085
rect 425 38275 595 38445
rect 425 38635 595 38805
rect 425 38995 595 39165
rect 425 39355 595 39525
rect 425 39715 595 39885
rect 65 31075 235 31245
rect 785 30715 955 30885
rect 785 31075 955 31245
rect 785 31435 955 31605
rect 785 31795 955 31965
rect 785 32155 955 32325
rect 785 32515 955 32685
rect 785 32875 955 33045
rect 785 33235 955 33405
rect 785 33595 955 33765
rect 785 33955 955 34125
rect 785 34315 955 34485
rect 785 34675 955 34845
rect 785 35035 955 35205
rect 785 35395 955 35565
rect 785 35755 955 35925
rect 785 36115 955 36285
rect 785 36475 955 36645
rect 785 36835 955 37005
rect 785 37195 955 37365
rect 785 37555 955 37725
rect 785 37915 955 38085
rect 785 38275 955 38445
rect 785 38635 955 38805
rect 785 38995 955 39165
rect 785 39355 955 39525
rect 785 39715 955 39885
rect 65 31435 235 31605
rect 65 31795 235 31965
rect 65 32155 235 32325
rect 1135 40280 1305 40450
rect 1495 40280 1665 40450
rect 1855 40280 2025 40450
rect 2215 40280 2385 40450
rect 2575 40280 2745 40450
rect 65 32515 235 32685
rect 65 32875 235 33045
rect 65 33235 235 33405
rect 65 33595 235 33765
rect 65 33955 235 34125
rect 65 34315 235 34485
rect 65 22435 235 22605
rect 65 22795 235 22965
rect 65 23155 235 23325
rect 65 23515 235 23685
rect 65 23875 235 24045
rect 65 20635 235 20805
rect 425 20635 595 20805
rect 425 20995 595 21165
rect 425 21355 595 21525
rect 425 21715 595 21885
rect 65 20995 235 21165
rect 785 20635 955 20805
rect 785 20995 955 21165
rect 785 21355 955 21525
rect 65 21715 235 21885
rect 785 21715 955 21885
rect 785 22075 955 22245
rect 785 22435 955 22605
rect 785 22795 955 22965
rect 785 23155 955 23325
rect 785 23515 955 23685
rect 785 23875 955 24045
rect 785 24235 955 24405
rect 785 24595 955 24765
rect 785 24955 955 25125
rect 785 25315 955 25485
rect 785 25675 955 25845
rect 785 26035 955 26205
rect 785 26395 955 26565
rect 785 26755 955 26925
rect 785 27115 955 27285
rect 785 27475 955 27645
rect 785 27835 955 28005
rect 785 28195 955 28365
rect 785 28555 955 28725
rect 785 28915 955 29085
rect 785 29275 955 29445
rect 785 29635 955 29805
rect 785 29995 955 30165
rect 425 22075 595 22245
rect 425 22435 595 22605
rect 425 22795 595 22965
rect 65 22075 235 22245
rect 425 23155 595 23325
rect 425 23515 595 23685
rect 425 23875 595 24045
rect 425 24235 595 24405
rect 425 24595 595 24765
rect 425 24955 595 25125
rect 425 25315 595 25485
rect 425 25675 595 25845
rect 425 26035 595 26205
rect 425 26395 595 26565
rect 425 26755 595 26925
rect 425 27115 595 27285
rect 425 27475 595 27645
rect 425 27835 595 28005
rect 425 28195 595 28365
rect 425 28555 595 28725
rect 425 28915 595 29085
rect 425 29275 595 29445
rect 425 29635 595 29805
rect 425 29995 595 30165
rect 65 24235 235 24405
rect 65 24595 235 24765
rect 65 24955 235 25125
rect 65 25315 235 25485
rect 65 21355 235 21525
rect 65 25675 235 25845
rect 65 26035 235 26205
rect 65 26395 235 26565
rect 65 26755 235 26925
rect 65 27115 235 27285
rect 65 27475 235 27645
rect 65 27835 235 28005
rect 65 28195 235 28365
rect 65 28555 235 28725
rect 65 28915 235 29085
rect 65 29275 235 29445
rect 65 29635 235 29805
rect 65 29995 235 30165
rect 5085 25315 5255 25485
rect 5085 25675 5255 25845
rect 5085 26035 5255 26205
rect 5085 26395 5255 26565
rect 5085 26755 5255 26925
rect 5085 27115 5255 27285
rect 5085 27475 5255 27645
rect 5085 27835 5255 28005
rect 5085 28195 5255 28365
rect 5085 28555 5255 28725
rect 5085 28915 5255 29085
rect 5085 29275 5255 29445
rect 5085 29635 5255 29805
rect 5085 29995 5255 30165
rect 5085 20635 5255 20805
rect 5445 20635 5615 20805
rect 5805 20635 5975 20805
rect 5805 20995 5975 21165
rect 5805 21355 5975 21525
rect 5805 21715 5975 21885
rect 5805 22075 5975 22245
rect 5805 22435 5975 22605
rect 5805 22795 5975 22965
rect 5805 23155 5975 23325
rect 5805 23515 5975 23685
rect 5805 23875 5975 24045
rect 5805 24235 5975 24405
rect 5805 24595 5975 24765
rect 5805 24955 5975 25125
rect 5805 25315 5975 25485
rect 5805 25675 5975 25845
rect 5805 26035 5975 26205
rect 5805 26395 5975 26565
rect 5805 26755 5975 26925
rect 5805 27115 5975 27285
rect 5805 27475 5975 27645
rect 5805 27835 5975 28005
rect 5805 28195 5975 28365
rect 5805 28555 5975 28725
rect 5805 28915 5975 29085
rect 5805 29275 5975 29445
rect 5805 29635 5975 29805
rect 5805 29995 5975 30165
rect 5445 20995 5615 21165
rect 5445 21355 5615 21525
rect 5445 21715 5615 21885
rect 5445 22075 5615 22245
rect 5445 22435 5615 22605
rect 5445 22795 5615 22965
rect 5445 23155 5615 23325
rect 5445 23515 5615 23685
rect 5445 23875 5615 24045
rect 5445 24235 5615 24405
rect 5445 24595 5615 24765
rect 5445 24955 5615 25125
rect 5445 25315 5615 25485
rect 5445 25675 5615 25845
rect 5445 26035 5615 26205
rect 5445 26395 5615 26565
rect 5445 26755 5615 26925
rect 5445 27115 5615 27285
rect 5445 27475 5615 27645
rect 5445 27835 5615 28005
rect 5445 28195 5615 28365
rect 5445 28555 5615 28725
rect 5445 28915 5615 29085
rect 5445 29275 5615 29445
rect 5445 29635 5615 29805
rect 5445 29995 5615 30165
rect 5085 20995 5255 21165
rect 5085 21355 5255 21525
rect 5085 21715 5255 21885
rect 5085 22075 5255 22245
rect 5085 22435 5255 22605
rect 5085 22795 5255 22965
rect 5085 23155 5255 23325
rect 5085 23515 5255 23685
rect 5085 23875 5255 24045
rect 5085 24235 5255 24405
rect 5085 24595 5255 24765
rect 5085 24955 5255 25125
rect 5085 10195 5255 10365
rect 65 10195 235 10365
rect 5445 10195 5615 10365
rect 785 10195 955 10365
rect 5805 10195 5975 10365
rect 425 10195 595 10365
rect 5085 12355 5255 12525
rect 5085 12715 5255 12885
rect 5085 13075 5255 13245
rect 5085 13435 5255 13605
rect 5085 13795 5255 13965
rect 5085 14155 5255 14325
rect 5085 14515 5255 14685
rect 5085 14875 5255 15045
rect 5085 15235 5255 15405
rect 5085 15595 5255 15765
rect 5085 15955 5255 16125
rect 5085 16315 5255 16485
rect 5085 16675 5255 16845
rect 5085 17035 5255 17205
rect 5085 17395 5255 17565
rect 5085 17755 5255 17925
rect 5085 18115 5255 18285
rect 5085 18475 5255 18645
rect 5085 18835 5255 19005
rect 5085 19195 5255 19365
rect 5085 19555 5255 19725
rect 5085 19915 5255 20085
rect 5085 10555 5255 10725
rect 5085 10915 5255 11085
rect 5445 10555 5615 10725
rect 5445 10915 5615 11085
rect 5445 11275 5615 11445
rect 5445 11635 5615 11805
rect 5445 11995 5615 12165
rect 5445 12355 5615 12525
rect 5445 12715 5615 12885
rect 5445 13075 5615 13245
rect 5445 13435 5615 13605
rect 5445 13795 5615 13965
rect 5445 14155 5615 14325
rect 5445 14515 5615 14685
rect 5445 14875 5615 15045
rect 5445 15235 5615 15405
rect 5445 15595 5615 15765
rect 5445 15955 5615 16125
rect 5445 16315 5615 16485
rect 5445 16675 5615 16845
rect 5445 17035 5615 17205
rect 5445 17395 5615 17565
rect 5445 17755 5615 17925
rect 5445 18115 5615 18285
rect 5445 18475 5615 18645
rect 5445 18835 5615 19005
rect 5445 19195 5615 19365
rect 5445 19555 5615 19725
rect 5445 19915 5615 20085
rect 5085 11275 5255 11445
rect 5085 11635 5255 11805
rect 5805 10555 5975 10725
rect 5805 10915 5975 11085
rect 5805 11275 5975 11445
rect 5805 11635 5975 11805
rect 5805 11995 5975 12165
rect 5805 12355 5975 12525
rect 5805 12715 5975 12885
rect 5805 13075 5975 13245
rect 5805 13435 5975 13605
rect 5805 13795 5975 13965
rect 5805 14155 5975 14325
rect 5805 14515 5975 14685
rect 5805 14875 5975 15045
rect 5805 15235 5975 15405
rect 5805 15595 5975 15765
rect 5805 15955 5975 16125
rect 5805 16315 5975 16485
rect 5805 16675 5975 16845
rect 5805 17035 5975 17205
rect 5805 17395 5975 17565
rect 5805 17755 5975 17925
rect 5805 18115 5975 18285
rect 5805 18475 5975 18645
rect 5805 18835 5975 19005
rect 5805 19195 5975 19365
rect 5805 19555 5975 19725
rect 5805 19915 5975 20085
rect 5085 11995 5255 12165
rect 785 10915 955 11085
rect 785 11275 955 11445
rect 785 11635 955 11805
rect 785 11995 955 12165
rect 785 12355 955 12525
rect 785 12715 955 12885
rect 785 13075 955 13245
rect 785 13435 955 13605
rect 785 13795 955 13965
rect 785 14155 955 14325
rect 785 14515 955 14685
rect 785 14875 955 15045
rect 785 15235 955 15405
rect 785 15595 955 15765
rect 785 15955 955 16125
rect 785 16315 955 16485
rect 785 16675 955 16845
rect 785 17035 955 17205
rect 785 17395 955 17565
rect 785 17755 955 17925
rect 785 18115 955 18285
rect 785 18475 955 18645
rect 785 18835 955 19005
rect 65 10555 235 10725
rect 65 10915 235 11085
rect 65 11275 235 11445
rect 65 11635 235 11805
rect 65 11995 235 12165
rect 65 12355 235 12525
rect 65 12715 235 12885
rect 65 13075 235 13245
rect 65 13435 235 13605
rect 65 13795 235 13965
rect 65 14155 235 14325
rect 65 14515 235 14685
rect 65 14875 235 15045
rect 65 15235 235 15405
rect 65 15595 235 15765
rect 65 15955 235 16125
rect 65 16315 235 16485
rect 65 16675 235 16845
rect 65 17035 235 17205
rect 65 17395 235 17565
rect 65 17755 235 17925
rect 65 18115 235 18285
rect 65 18475 235 18645
rect 425 19915 595 20085
rect 65 19915 235 20085
rect 65 18835 235 19005
rect 65 19195 235 19365
rect 425 19555 595 19725
rect 785 19195 955 19365
rect 785 19555 955 19725
rect 785 19915 955 20085
rect 65 19555 235 19725
rect 785 10555 955 10725
rect 425 10555 595 10725
rect 425 10915 595 11085
rect 425 11275 595 11445
rect 425 11635 595 11805
rect 425 11995 595 12165
rect 425 12355 595 12525
rect 425 12715 595 12885
rect 425 13075 595 13245
rect 425 13435 595 13605
rect 425 13795 595 13965
rect 425 14155 595 14325
rect 425 14515 595 14685
rect 425 14875 595 15045
rect 425 15235 595 15405
rect 425 15595 595 15765
rect 425 15955 595 16125
rect 425 16315 595 16485
rect 425 16675 595 16845
rect 425 17035 595 17205
rect 425 17395 595 17565
rect 425 17755 595 17925
rect 425 18115 595 18285
rect 425 18475 595 18645
rect 425 18835 595 19005
rect 425 19195 595 19365
rect 65 9115 235 9285
rect 785 115 955 285
rect 785 475 955 645
rect 785 835 955 1005
rect 785 1195 955 1365
rect 785 1555 955 1725
rect 785 1915 955 2085
rect 785 2275 955 2445
rect 785 2635 955 2805
rect 785 2995 955 3165
rect 785 3355 955 3525
rect 785 3715 955 3885
rect 785 4075 955 4245
rect 785 4435 955 4605
rect 785 4795 955 4965
rect 785 5155 955 5325
rect 785 5515 955 5685
rect 785 5875 955 6045
rect 785 6235 955 6405
rect 785 6595 955 6765
rect 785 6955 955 7125
rect 785 7315 955 7485
rect 785 7675 955 7845
rect 785 8035 955 8205
rect 785 8395 955 8565
rect 785 8755 955 8925
rect 785 9115 955 9285
rect 785 9475 955 9645
rect 785 9835 955 10005
rect 65 9475 235 9645
rect 425 115 595 285
rect 425 475 595 645
rect 425 835 595 1005
rect 425 1195 595 1365
rect 425 1555 595 1725
rect 425 1915 595 2085
rect 425 2275 595 2445
rect 425 2635 595 2805
rect 425 2995 595 3165
rect 425 3355 595 3525
rect 425 3715 595 3885
rect 425 4075 595 4245
rect 425 4435 595 4605
rect 425 4795 595 4965
rect 425 5155 595 5325
rect 425 5515 595 5685
rect 425 5875 595 6045
rect 425 6235 595 6405
rect 425 6595 595 6765
rect 425 6955 595 7125
rect 425 7315 595 7485
rect 425 7675 595 7845
rect 425 8035 595 8205
rect 425 8395 595 8565
rect 425 8755 595 8925
rect 425 9115 595 9285
rect 425 9475 595 9645
rect 425 9835 595 10005
rect 65 9835 235 10005
rect 65 115 235 285
rect 65 475 235 645
rect 65 835 235 1005
rect 65 1195 235 1365
rect 65 1555 235 1725
rect 65 1915 235 2085
rect 65 2275 235 2445
rect 65 2635 235 2805
rect 65 2995 235 3165
rect 65 3355 235 3525
rect 65 3715 235 3885
rect 65 4075 235 4245
rect 65 4435 235 4605
rect 65 4795 235 4965
rect 65 5155 235 5325
rect 65 5515 235 5685
rect 65 5875 235 6045
rect 65 6235 235 6405
rect 65 6595 235 6765
rect 65 6955 235 7125
rect 65 7315 235 7485
rect 65 7675 235 7845
rect 65 8035 235 8205
rect 65 8395 235 8565
rect 65 8755 235 8925
rect 5445 9115 5615 9285
rect 5445 9475 5615 9645
rect 5445 9835 5615 10005
rect 5085 4075 5255 4245
rect 5085 4435 5255 4605
rect 5085 4795 5255 4965
rect 5085 5155 5255 5325
rect 5085 5515 5255 5685
rect 5085 5875 5255 6045
rect 5085 6235 5255 6405
rect 5085 6595 5255 6765
rect 5085 6955 5255 7125
rect 5085 7315 5255 7485
rect 5085 7675 5255 7845
rect 5085 8035 5255 8205
rect 5085 8395 5255 8565
rect 5085 8755 5255 8925
rect 5085 9115 5255 9285
rect 5085 9475 5255 9645
rect 5085 9835 5255 10005
rect 5085 2995 5255 3165
rect 5085 3355 5255 3525
rect 5085 3715 5255 3885
rect 5445 115 5615 285
rect 5445 475 5615 645
rect 5445 835 5615 1005
rect 5445 1195 5615 1365
rect 5445 1555 5615 1725
rect 5445 1915 5615 2085
rect 5445 2275 5615 2445
rect 5445 2635 5615 2805
rect 5445 2995 5615 3165
rect 5445 3355 5615 3525
rect 5445 3715 5615 3885
rect 5445 4075 5615 4245
rect 5445 4435 5615 4605
rect 5445 4795 5615 4965
rect 5445 5155 5615 5325
rect 5805 115 5975 285
rect 5805 475 5975 645
rect 5805 835 5975 1005
rect 5805 1195 5975 1365
rect 5805 1555 5975 1725
rect 5805 1915 5975 2085
rect 5805 2275 5975 2445
rect 5805 2635 5975 2805
rect 5805 2995 5975 3165
rect 5805 3355 5975 3525
rect 5805 3715 5975 3885
rect 5805 4075 5975 4245
rect 5805 4435 5975 4605
rect 5805 4795 5975 4965
rect 5805 5155 5975 5325
rect 5805 5515 5975 5685
rect 5805 5875 5975 6045
rect 5805 6235 5975 6405
rect 5805 6595 5975 6765
rect 5805 6955 5975 7125
rect 5805 7315 5975 7485
rect 5805 7675 5975 7845
rect 5805 8035 5975 8205
rect 5805 8395 5975 8565
rect 5805 8755 5975 8925
rect 5805 9115 5975 9285
rect 5805 9475 5975 9645
rect 5805 9835 5975 10005
rect 5445 5515 5615 5685
rect 5445 5875 5615 6045
rect 5445 6235 5615 6405
rect 5445 6595 5615 6765
rect 5445 6955 5615 7125
rect 5445 7315 5615 7485
rect 5445 7675 5615 7845
rect 5445 8035 5615 8205
rect 5445 8395 5615 8565
rect 5445 8755 5615 8925
rect 5085 115 5255 285
rect 5085 475 5255 645
rect 5085 835 5255 1005
rect 5085 1195 5255 1365
rect 5085 1555 5255 1725
rect 5085 1915 5255 2085
rect 5085 2275 5255 2445
rect 5085 2635 5255 2805
<< l95d20 >>
rect 1010 40190 5030 40540
<< l67d20 >>
rect 65 35 955 39965
rect 5085 35 5975 39965
rect 1055 40280 4985 40450
rect 6258 35 7148 39965
<< l68d20 >>
rect 35 55 985 39945
rect 5055 55 6005 39945
rect 1075 40250 4965 40480
<< l65d20 >>
rect 0 0 6040 40000
<< l93d44 >>
rect 6040 -125 7492 40125
<< l64d20 >>
rect -305 -380 7671 40720
<< l65d44 >>
rect 6040 0 7366 40000
<< end >>
