magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< error_s >>
rect 97 996 6233 1039
rect 165 307 403 329
<< viali >>
rect 188 2309 8142 2487
rect 196 53 230 87
rect 268 53 302 87
<< metal1 >>
rect 172 2444 179 2496
rect 231 2487 251 2496
rect 303 2487 323 2496
rect 375 2487 395 2496
rect 447 2487 467 2496
rect 519 2487 539 2496
rect 591 2487 611 2496
rect 663 2487 683 2496
rect 735 2487 755 2496
rect 807 2487 827 2496
rect 879 2487 899 2496
rect 951 2487 971 2496
rect 1023 2487 1043 2496
rect 1095 2487 1115 2496
rect 1167 2487 1187 2496
rect 1239 2487 1259 2496
rect 1311 2487 1331 2496
rect 1383 2487 1403 2496
rect 1455 2487 1475 2496
rect 1527 2487 1547 2496
rect 1599 2487 1619 2496
rect 1671 2487 1691 2496
rect 1743 2487 1763 2496
rect 1815 2487 1835 2496
rect 1887 2487 1907 2496
rect 1959 2487 1979 2496
rect 2031 2487 2051 2496
rect 2103 2487 2123 2496
rect 2175 2487 2195 2496
rect 2247 2487 2267 2496
rect 2319 2487 2339 2496
rect 2391 2487 2411 2496
rect 2463 2487 2483 2496
rect 2535 2487 2555 2496
rect 2607 2487 2627 2496
rect 2679 2487 2699 2496
rect 2751 2487 2771 2496
rect 2823 2487 2843 2496
rect 2895 2487 2915 2496
rect 2967 2487 2987 2496
rect 3039 2487 3059 2496
rect 3111 2487 3131 2496
rect 3183 2487 3203 2496
rect 3255 2487 3275 2496
rect 3327 2487 3347 2496
rect 3399 2487 3419 2496
rect 3471 2487 3491 2496
rect 3543 2487 3563 2496
rect 3615 2487 3635 2496
rect 3687 2487 3707 2496
rect 3759 2487 3779 2496
rect 3831 2487 3851 2496
rect 3903 2487 3923 2496
rect 3975 2487 3995 2496
rect 4047 2487 4067 2496
rect 4119 2487 4139 2496
rect 4191 2487 4211 2496
rect 4263 2487 4283 2496
rect 4335 2487 4355 2496
rect 4407 2487 4427 2496
rect 4479 2487 4499 2496
rect 4551 2487 4571 2496
rect 4623 2487 4643 2496
rect 4695 2487 4715 2496
rect 4767 2487 4787 2496
rect 4839 2487 4859 2496
rect 4911 2487 4931 2496
rect 4983 2487 5003 2496
rect 5055 2487 5075 2496
rect 5127 2487 5147 2496
rect 5199 2487 5219 2496
rect 5271 2487 5291 2496
rect 5343 2487 5363 2496
rect 5415 2487 5435 2496
rect 5487 2487 5507 2496
rect 5559 2487 5579 2496
rect 5631 2487 5651 2496
rect 5703 2487 5723 2496
rect 5775 2487 5795 2496
rect 5847 2487 5867 2496
rect 5919 2487 5939 2496
rect 5991 2487 6011 2496
rect 6063 2487 6083 2496
rect 6135 2487 6155 2496
rect 6207 2487 6227 2496
rect 6279 2487 6299 2496
rect 6351 2487 6371 2496
rect 6423 2487 6443 2496
rect 6495 2487 6515 2496
rect 6567 2487 6587 2496
rect 6639 2487 6659 2496
rect 6711 2487 6731 2496
rect 6783 2487 6803 2496
rect 6855 2487 6875 2496
rect 6927 2487 6947 2496
rect 6999 2487 7019 2496
rect 7071 2487 7091 2496
rect 7143 2487 7163 2496
rect 7215 2487 7235 2496
rect 7287 2487 7307 2496
rect 7359 2487 7379 2496
rect 7431 2487 7451 2496
rect 7503 2487 7523 2496
rect 7575 2487 7595 2496
rect 7647 2487 7667 2496
rect 7719 2487 7739 2496
rect 7791 2487 7811 2496
rect 7863 2487 7883 2496
rect 7935 2487 7955 2496
rect 8007 2487 8027 2496
rect 8079 2487 8099 2496
rect 8151 2444 8158 2496
rect 172 2424 188 2444
rect 8142 2424 8158 2444
rect 172 2372 179 2424
rect 8151 2372 8158 2424
rect 172 2352 188 2372
rect 8142 2352 8158 2372
rect 172 2309 179 2352
rect 8151 2309 8158 2352
rect 176 2300 179 2309
rect 231 2300 251 2309
rect 303 2300 323 2309
rect 375 2300 395 2309
rect 447 2300 467 2309
rect 519 2300 539 2309
rect 591 2300 611 2309
rect 663 2300 683 2309
rect 735 2300 755 2309
rect 807 2300 827 2309
rect 879 2300 899 2309
rect 951 2300 971 2309
rect 1023 2300 1043 2309
rect 1095 2300 1115 2309
rect 1167 2300 1187 2309
rect 1239 2300 1259 2309
rect 1311 2300 1331 2309
rect 1383 2300 1403 2309
rect 1455 2300 1475 2309
rect 1527 2300 1547 2309
rect 1599 2300 1619 2309
rect 1671 2300 1691 2309
rect 1743 2300 1763 2309
rect 1815 2300 1835 2309
rect 1887 2300 1907 2309
rect 1959 2300 1979 2309
rect 2031 2300 2051 2309
rect 2103 2300 2123 2309
rect 2175 2300 2195 2309
rect 2247 2300 2267 2309
rect 2319 2300 2339 2309
rect 2391 2300 2411 2309
rect 2463 2300 2483 2309
rect 2535 2300 2555 2309
rect 2607 2300 2627 2309
rect 2679 2300 2699 2309
rect 2751 2300 2771 2309
rect 2823 2300 2843 2309
rect 2895 2300 2915 2309
rect 2967 2300 2987 2309
rect 3039 2300 3059 2309
rect 3111 2300 3131 2309
rect 3183 2300 3203 2309
rect 3255 2300 3275 2309
rect 3327 2300 3347 2309
rect 3399 2300 3419 2309
rect 3471 2300 3491 2309
rect 3543 2300 3563 2309
rect 3615 2300 3635 2309
rect 3687 2300 3707 2309
rect 3759 2300 3779 2309
rect 3831 2300 3851 2309
rect 3903 2300 3923 2309
rect 3975 2300 3995 2309
rect 4047 2300 4067 2309
rect 4119 2300 4139 2309
rect 4191 2300 4211 2309
rect 4263 2300 4283 2309
rect 4335 2300 4355 2309
rect 4407 2300 4427 2309
rect 4479 2300 4499 2309
rect 4551 2300 4571 2309
rect 4623 2300 4643 2309
rect 4695 2300 4715 2309
rect 4767 2300 4787 2309
rect 4839 2300 4859 2309
rect 4911 2300 4931 2309
rect 4983 2300 5003 2309
rect 5055 2300 5075 2309
rect 5127 2300 5147 2309
rect 5199 2300 5219 2309
rect 5271 2300 5291 2309
rect 5343 2300 5363 2309
rect 5415 2300 5435 2309
rect 5487 2300 5507 2309
rect 5559 2300 5579 2309
rect 5631 2300 5651 2309
rect 5703 2300 5723 2309
rect 5775 2300 5795 2309
rect 5847 2300 5867 2309
rect 5919 2300 5939 2309
rect 5991 2300 6011 2309
rect 6063 2300 6083 2309
rect 6135 2300 6155 2309
rect 6207 2300 6227 2309
rect 6279 2300 6299 2309
rect 6351 2300 6371 2309
rect 6423 2300 6443 2309
rect 6495 2300 6515 2309
rect 6567 2300 6587 2309
rect 6639 2300 6659 2309
rect 6711 2300 6731 2309
rect 6783 2300 6803 2309
rect 6855 2300 6875 2309
rect 6927 2300 6947 2309
rect 6999 2300 7019 2309
rect 7071 2300 7091 2309
rect 7143 2300 7163 2309
rect 7215 2300 7235 2309
rect 7287 2300 7307 2309
rect 7359 2300 7379 2309
rect 7431 2300 7451 2309
rect 7503 2300 7523 2309
rect 7575 2300 7595 2309
rect 7647 2300 7667 2309
rect 7719 2300 7739 2309
rect 7791 2300 7811 2309
rect 7863 2300 7883 2309
rect 7935 2300 7955 2309
rect 8007 2300 8027 2309
rect 8079 2300 8099 2309
rect 8151 2300 8154 2309
rect 176 2258 8154 2300
rect 0 466 115 2050
rect 176 846 8154 1254
rect 8 127 144 263
rect 180 222 318 432
rect 180 162 318 168
rect 180 110 186 162
rect 238 110 260 162
rect 312 110 318 162
rect 180 88 318 110
rect 180 36 186 88
rect 238 36 260 88
rect 312 36 318 88
rect 180 30 318 36
<< via1 >>
rect 179 2487 231 2496
rect 251 2487 303 2496
rect 323 2487 375 2496
rect 395 2487 447 2496
rect 467 2487 519 2496
rect 539 2487 591 2496
rect 611 2487 663 2496
rect 683 2487 735 2496
rect 755 2487 807 2496
rect 827 2487 879 2496
rect 899 2487 951 2496
rect 971 2487 1023 2496
rect 1043 2487 1095 2496
rect 1115 2487 1167 2496
rect 1187 2487 1239 2496
rect 1259 2487 1311 2496
rect 1331 2487 1383 2496
rect 1403 2487 1455 2496
rect 1475 2487 1527 2496
rect 1547 2487 1599 2496
rect 1619 2487 1671 2496
rect 1691 2487 1743 2496
rect 1763 2487 1815 2496
rect 1835 2487 1887 2496
rect 1907 2487 1959 2496
rect 1979 2487 2031 2496
rect 2051 2487 2103 2496
rect 2123 2487 2175 2496
rect 2195 2487 2247 2496
rect 2267 2487 2319 2496
rect 2339 2487 2391 2496
rect 2411 2487 2463 2496
rect 2483 2487 2535 2496
rect 2555 2487 2607 2496
rect 2627 2487 2679 2496
rect 2699 2487 2751 2496
rect 2771 2487 2823 2496
rect 2843 2487 2895 2496
rect 2915 2487 2967 2496
rect 2987 2487 3039 2496
rect 3059 2487 3111 2496
rect 3131 2487 3183 2496
rect 3203 2487 3255 2496
rect 3275 2487 3327 2496
rect 3347 2487 3399 2496
rect 3419 2487 3471 2496
rect 3491 2487 3543 2496
rect 3563 2487 3615 2496
rect 3635 2487 3687 2496
rect 3707 2487 3759 2496
rect 3779 2487 3831 2496
rect 3851 2487 3903 2496
rect 3923 2487 3975 2496
rect 3995 2487 4047 2496
rect 4067 2487 4119 2496
rect 4139 2487 4191 2496
rect 4211 2487 4263 2496
rect 4283 2487 4335 2496
rect 4355 2487 4407 2496
rect 4427 2487 4479 2496
rect 4499 2487 4551 2496
rect 4571 2487 4623 2496
rect 4643 2487 4695 2496
rect 4715 2487 4767 2496
rect 4787 2487 4839 2496
rect 4859 2487 4911 2496
rect 4931 2487 4983 2496
rect 5003 2487 5055 2496
rect 5075 2487 5127 2496
rect 5147 2487 5199 2496
rect 5219 2487 5271 2496
rect 5291 2487 5343 2496
rect 5363 2487 5415 2496
rect 5435 2487 5487 2496
rect 5507 2487 5559 2496
rect 5579 2487 5631 2496
rect 5651 2487 5703 2496
rect 5723 2487 5775 2496
rect 5795 2487 5847 2496
rect 5867 2487 5919 2496
rect 5939 2487 5991 2496
rect 6011 2487 6063 2496
rect 6083 2487 6135 2496
rect 6155 2487 6207 2496
rect 6227 2487 6279 2496
rect 6299 2487 6351 2496
rect 6371 2487 6423 2496
rect 6443 2487 6495 2496
rect 6515 2487 6567 2496
rect 6587 2487 6639 2496
rect 6659 2487 6711 2496
rect 6731 2487 6783 2496
rect 6803 2487 6855 2496
rect 6875 2487 6927 2496
rect 6947 2487 6999 2496
rect 7019 2487 7071 2496
rect 7091 2487 7143 2496
rect 7163 2487 7215 2496
rect 7235 2487 7287 2496
rect 7307 2487 7359 2496
rect 7379 2487 7431 2496
rect 7451 2487 7503 2496
rect 7523 2487 7575 2496
rect 7595 2487 7647 2496
rect 7667 2487 7719 2496
rect 7739 2487 7791 2496
rect 7811 2487 7863 2496
rect 7883 2487 7935 2496
rect 7955 2487 8007 2496
rect 8027 2487 8079 2496
rect 8099 2487 8151 2496
rect 179 2444 188 2487
rect 188 2444 231 2487
rect 251 2444 303 2487
rect 323 2444 375 2487
rect 395 2444 447 2487
rect 467 2444 519 2487
rect 539 2444 591 2487
rect 611 2444 663 2487
rect 683 2444 735 2487
rect 755 2444 807 2487
rect 827 2444 879 2487
rect 899 2444 951 2487
rect 971 2444 1023 2487
rect 1043 2444 1095 2487
rect 1115 2444 1167 2487
rect 1187 2444 1239 2487
rect 1259 2444 1311 2487
rect 1331 2444 1383 2487
rect 1403 2444 1455 2487
rect 1475 2444 1527 2487
rect 1547 2444 1599 2487
rect 1619 2444 1671 2487
rect 1691 2444 1743 2487
rect 1763 2444 1815 2487
rect 1835 2444 1887 2487
rect 1907 2444 1959 2487
rect 1979 2444 2031 2487
rect 2051 2444 2103 2487
rect 2123 2444 2175 2487
rect 2195 2444 2247 2487
rect 2267 2444 2319 2487
rect 2339 2444 2391 2487
rect 2411 2444 2463 2487
rect 2483 2444 2535 2487
rect 2555 2444 2607 2487
rect 2627 2444 2679 2487
rect 2699 2444 2751 2487
rect 2771 2444 2823 2487
rect 2843 2444 2895 2487
rect 2915 2444 2967 2487
rect 2987 2444 3039 2487
rect 3059 2444 3111 2487
rect 3131 2444 3183 2487
rect 3203 2444 3255 2487
rect 3275 2444 3327 2487
rect 3347 2444 3399 2487
rect 3419 2444 3471 2487
rect 3491 2444 3543 2487
rect 3563 2444 3615 2487
rect 3635 2444 3687 2487
rect 3707 2444 3759 2487
rect 3779 2444 3831 2487
rect 3851 2444 3903 2487
rect 3923 2444 3975 2487
rect 3995 2444 4047 2487
rect 4067 2444 4119 2487
rect 4139 2444 4191 2487
rect 4211 2444 4263 2487
rect 4283 2444 4335 2487
rect 4355 2444 4407 2487
rect 4427 2444 4479 2487
rect 4499 2444 4551 2487
rect 4571 2444 4623 2487
rect 4643 2444 4695 2487
rect 4715 2444 4767 2487
rect 4787 2444 4839 2487
rect 4859 2444 4911 2487
rect 4931 2444 4983 2487
rect 5003 2444 5055 2487
rect 5075 2444 5127 2487
rect 5147 2444 5199 2487
rect 5219 2444 5271 2487
rect 5291 2444 5343 2487
rect 5363 2444 5415 2487
rect 5435 2444 5487 2487
rect 5507 2444 5559 2487
rect 5579 2444 5631 2487
rect 5651 2444 5703 2487
rect 5723 2444 5775 2487
rect 5795 2444 5847 2487
rect 5867 2444 5919 2487
rect 5939 2444 5991 2487
rect 6011 2444 6063 2487
rect 6083 2444 6135 2487
rect 6155 2444 6207 2487
rect 6227 2444 6279 2487
rect 6299 2444 6351 2487
rect 6371 2444 6423 2487
rect 6443 2444 6495 2487
rect 6515 2444 6567 2487
rect 6587 2444 6639 2487
rect 6659 2444 6711 2487
rect 6731 2444 6783 2487
rect 6803 2444 6855 2487
rect 6875 2444 6927 2487
rect 6947 2444 6999 2487
rect 7019 2444 7071 2487
rect 7091 2444 7143 2487
rect 7163 2444 7215 2487
rect 7235 2444 7287 2487
rect 7307 2444 7359 2487
rect 7379 2444 7431 2487
rect 7451 2444 7503 2487
rect 7523 2444 7575 2487
rect 7595 2444 7647 2487
rect 7667 2444 7719 2487
rect 7739 2444 7791 2487
rect 7811 2444 7863 2487
rect 7883 2444 7935 2487
rect 7955 2444 8007 2487
rect 8027 2444 8079 2487
rect 8099 2444 8142 2487
rect 8142 2444 8151 2487
rect 179 2372 188 2424
rect 188 2372 231 2424
rect 251 2372 303 2424
rect 323 2372 375 2424
rect 395 2372 447 2424
rect 467 2372 519 2424
rect 539 2372 591 2424
rect 611 2372 663 2424
rect 683 2372 735 2424
rect 755 2372 807 2424
rect 827 2372 879 2424
rect 899 2372 951 2424
rect 971 2372 1023 2424
rect 1043 2372 1095 2424
rect 1115 2372 1167 2424
rect 1187 2372 1239 2424
rect 1259 2372 1311 2424
rect 1331 2372 1383 2424
rect 1403 2372 1455 2424
rect 1475 2372 1527 2424
rect 1547 2372 1599 2424
rect 1619 2372 1671 2424
rect 1691 2372 1743 2424
rect 1763 2372 1815 2424
rect 1835 2372 1887 2424
rect 1907 2372 1959 2424
rect 1979 2372 2031 2424
rect 2051 2372 2103 2424
rect 2123 2372 2175 2424
rect 2195 2372 2247 2424
rect 2267 2372 2319 2424
rect 2339 2372 2391 2424
rect 2411 2372 2463 2424
rect 2483 2372 2535 2424
rect 2555 2372 2607 2424
rect 2627 2372 2679 2424
rect 2699 2372 2751 2424
rect 2771 2372 2823 2424
rect 2843 2372 2895 2424
rect 2915 2372 2967 2424
rect 2987 2372 3039 2424
rect 3059 2372 3111 2424
rect 3131 2372 3183 2424
rect 3203 2372 3255 2424
rect 3275 2372 3327 2424
rect 3347 2372 3399 2424
rect 3419 2372 3471 2424
rect 3491 2372 3543 2424
rect 3563 2372 3615 2424
rect 3635 2372 3687 2424
rect 3707 2372 3759 2424
rect 3779 2372 3831 2424
rect 3851 2372 3903 2424
rect 3923 2372 3975 2424
rect 3995 2372 4047 2424
rect 4067 2372 4119 2424
rect 4139 2372 4191 2424
rect 4211 2372 4263 2424
rect 4283 2372 4335 2424
rect 4355 2372 4407 2424
rect 4427 2372 4479 2424
rect 4499 2372 4551 2424
rect 4571 2372 4623 2424
rect 4643 2372 4695 2424
rect 4715 2372 4767 2424
rect 4787 2372 4839 2424
rect 4859 2372 4911 2424
rect 4931 2372 4983 2424
rect 5003 2372 5055 2424
rect 5075 2372 5127 2424
rect 5147 2372 5199 2424
rect 5219 2372 5271 2424
rect 5291 2372 5343 2424
rect 5363 2372 5415 2424
rect 5435 2372 5487 2424
rect 5507 2372 5559 2424
rect 5579 2372 5631 2424
rect 5651 2372 5703 2424
rect 5723 2372 5775 2424
rect 5795 2372 5847 2424
rect 5867 2372 5919 2424
rect 5939 2372 5991 2424
rect 6011 2372 6063 2424
rect 6083 2372 6135 2424
rect 6155 2372 6207 2424
rect 6227 2372 6279 2424
rect 6299 2372 6351 2424
rect 6371 2372 6423 2424
rect 6443 2372 6495 2424
rect 6515 2372 6567 2424
rect 6587 2372 6639 2424
rect 6659 2372 6711 2424
rect 6731 2372 6783 2424
rect 6803 2372 6855 2424
rect 6875 2372 6927 2424
rect 6947 2372 6999 2424
rect 7019 2372 7071 2424
rect 7091 2372 7143 2424
rect 7163 2372 7215 2424
rect 7235 2372 7287 2424
rect 7307 2372 7359 2424
rect 7379 2372 7431 2424
rect 7451 2372 7503 2424
rect 7523 2372 7575 2424
rect 7595 2372 7647 2424
rect 7667 2372 7719 2424
rect 7739 2372 7791 2424
rect 7811 2372 7863 2424
rect 7883 2372 7935 2424
rect 7955 2372 8007 2424
rect 8027 2372 8079 2424
rect 8099 2372 8142 2424
rect 8142 2372 8151 2424
rect 179 2309 188 2352
rect 188 2309 231 2352
rect 251 2309 303 2352
rect 323 2309 375 2352
rect 395 2309 447 2352
rect 467 2309 519 2352
rect 539 2309 591 2352
rect 611 2309 663 2352
rect 683 2309 735 2352
rect 755 2309 807 2352
rect 827 2309 879 2352
rect 899 2309 951 2352
rect 971 2309 1023 2352
rect 1043 2309 1095 2352
rect 1115 2309 1167 2352
rect 1187 2309 1239 2352
rect 1259 2309 1311 2352
rect 1331 2309 1383 2352
rect 1403 2309 1455 2352
rect 1475 2309 1527 2352
rect 1547 2309 1599 2352
rect 1619 2309 1671 2352
rect 1691 2309 1743 2352
rect 1763 2309 1815 2352
rect 1835 2309 1887 2352
rect 1907 2309 1959 2352
rect 1979 2309 2031 2352
rect 2051 2309 2103 2352
rect 2123 2309 2175 2352
rect 2195 2309 2247 2352
rect 2267 2309 2319 2352
rect 2339 2309 2391 2352
rect 2411 2309 2463 2352
rect 2483 2309 2535 2352
rect 2555 2309 2607 2352
rect 2627 2309 2679 2352
rect 2699 2309 2751 2352
rect 2771 2309 2823 2352
rect 2843 2309 2895 2352
rect 2915 2309 2967 2352
rect 2987 2309 3039 2352
rect 3059 2309 3111 2352
rect 3131 2309 3183 2352
rect 3203 2309 3255 2352
rect 3275 2309 3327 2352
rect 3347 2309 3399 2352
rect 3419 2309 3471 2352
rect 3491 2309 3543 2352
rect 3563 2309 3615 2352
rect 3635 2309 3687 2352
rect 3707 2309 3759 2352
rect 3779 2309 3831 2352
rect 3851 2309 3903 2352
rect 3923 2309 3975 2352
rect 3995 2309 4047 2352
rect 4067 2309 4119 2352
rect 4139 2309 4191 2352
rect 4211 2309 4263 2352
rect 4283 2309 4335 2352
rect 4355 2309 4407 2352
rect 4427 2309 4479 2352
rect 4499 2309 4551 2352
rect 4571 2309 4623 2352
rect 4643 2309 4695 2352
rect 4715 2309 4767 2352
rect 4787 2309 4839 2352
rect 4859 2309 4911 2352
rect 4931 2309 4983 2352
rect 5003 2309 5055 2352
rect 5075 2309 5127 2352
rect 5147 2309 5199 2352
rect 5219 2309 5271 2352
rect 5291 2309 5343 2352
rect 5363 2309 5415 2352
rect 5435 2309 5487 2352
rect 5507 2309 5559 2352
rect 5579 2309 5631 2352
rect 5651 2309 5703 2352
rect 5723 2309 5775 2352
rect 5795 2309 5847 2352
rect 5867 2309 5919 2352
rect 5939 2309 5991 2352
rect 6011 2309 6063 2352
rect 6083 2309 6135 2352
rect 6155 2309 6207 2352
rect 6227 2309 6279 2352
rect 6299 2309 6351 2352
rect 6371 2309 6423 2352
rect 6443 2309 6495 2352
rect 6515 2309 6567 2352
rect 6587 2309 6639 2352
rect 6659 2309 6711 2352
rect 6731 2309 6783 2352
rect 6803 2309 6855 2352
rect 6875 2309 6927 2352
rect 6947 2309 6999 2352
rect 7019 2309 7071 2352
rect 7091 2309 7143 2352
rect 7163 2309 7215 2352
rect 7235 2309 7287 2352
rect 7307 2309 7359 2352
rect 7379 2309 7431 2352
rect 7451 2309 7503 2352
rect 7523 2309 7575 2352
rect 7595 2309 7647 2352
rect 7667 2309 7719 2352
rect 7739 2309 7791 2352
rect 7811 2309 7863 2352
rect 7883 2309 7935 2352
rect 7955 2309 8007 2352
rect 8027 2309 8079 2352
rect 8099 2309 8142 2352
rect 8142 2309 8151 2352
rect 179 2300 231 2309
rect 251 2300 303 2309
rect 323 2300 375 2309
rect 395 2300 447 2309
rect 467 2300 519 2309
rect 539 2300 591 2309
rect 611 2300 663 2309
rect 683 2300 735 2309
rect 755 2300 807 2309
rect 827 2300 879 2309
rect 899 2300 951 2309
rect 971 2300 1023 2309
rect 1043 2300 1095 2309
rect 1115 2300 1167 2309
rect 1187 2300 1239 2309
rect 1259 2300 1311 2309
rect 1331 2300 1383 2309
rect 1403 2300 1455 2309
rect 1475 2300 1527 2309
rect 1547 2300 1599 2309
rect 1619 2300 1671 2309
rect 1691 2300 1743 2309
rect 1763 2300 1815 2309
rect 1835 2300 1887 2309
rect 1907 2300 1959 2309
rect 1979 2300 2031 2309
rect 2051 2300 2103 2309
rect 2123 2300 2175 2309
rect 2195 2300 2247 2309
rect 2267 2300 2319 2309
rect 2339 2300 2391 2309
rect 2411 2300 2463 2309
rect 2483 2300 2535 2309
rect 2555 2300 2607 2309
rect 2627 2300 2679 2309
rect 2699 2300 2751 2309
rect 2771 2300 2823 2309
rect 2843 2300 2895 2309
rect 2915 2300 2967 2309
rect 2987 2300 3039 2309
rect 3059 2300 3111 2309
rect 3131 2300 3183 2309
rect 3203 2300 3255 2309
rect 3275 2300 3327 2309
rect 3347 2300 3399 2309
rect 3419 2300 3471 2309
rect 3491 2300 3543 2309
rect 3563 2300 3615 2309
rect 3635 2300 3687 2309
rect 3707 2300 3759 2309
rect 3779 2300 3831 2309
rect 3851 2300 3903 2309
rect 3923 2300 3975 2309
rect 3995 2300 4047 2309
rect 4067 2300 4119 2309
rect 4139 2300 4191 2309
rect 4211 2300 4263 2309
rect 4283 2300 4335 2309
rect 4355 2300 4407 2309
rect 4427 2300 4479 2309
rect 4499 2300 4551 2309
rect 4571 2300 4623 2309
rect 4643 2300 4695 2309
rect 4715 2300 4767 2309
rect 4787 2300 4839 2309
rect 4859 2300 4911 2309
rect 4931 2300 4983 2309
rect 5003 2300 5055 2309
rect 5075 2300 5127 2309
rect 5147 2300 5199 2309
rect 5219 2300 5271 2309
rect 5291 2300 5343 2309
rect 5363 2300 5415 2309
rect 5435 2300 5487 2309
rect 5507 2300 5559 2309
rect 5579 2300 5631 2309
rect 5651 2300 5703 2309
rect 5723 2300 5775 2309
rect 5795 2300 5847 2309
rect 5867 2300 5919 2309
rect 5939 2300 5991 2309
rect 6011 2300 6063 2309
rect 6083 2300 6135 2309
rect 6155 2300 6207 2309
rect 6227 2300 6279 2309
rect 6299 2300 6351 2309
rect 6371 2300 6423 2309
rect 6443 2300 6495 2309
rect 6515 2300 6567 2309
rect 6587 2300 6639 2309
rect 6659 2300 6711 2309
rect 6731 2300 6783 2309
rect 6803 2300 6855 2309
rect 6875 2300 6927 2309
rect 6947 2300 6999 2309
rect 7019 2300 7071 2309
rect 7091 2300 7143 2309
rect 7163 2300 7215 2309
rect 7235 2300 7287 2309
rect 7307 2300 7359 2309
rect 7379 2300 7431 2309
rect 7451 2300 7503 2309
rect 7523 2300 7575 2309
rect 7595 2300 7647 2309
rect 7667 2300 7719 2309
rect 7739 2300 7791 2309
rect 7811 2300 7863 2309
rect 7883 2300 7935 2309
rect 7955 2300 8007 2309
rect 8027 2300 8079 2309
rect 8099 2300 8151 2309
rect 186 110 238 162
rect 260 110 312 162
rect 186 87 238 88
rect 186 53 196 87
rect 196 53 230 87
rect 230 53 238 87
rect 186 36 238 53
rect 260 87 312 88
rect 260 53 268 87
rect 268 53 302 87
rect 302 53 312 87
rect 260 36 312 53
<< metal2 >>
rect 173 2496 8157 2502
rect 173 2444 179 2496
rect 231 2444 251 2496
rect 303 2444 323 2496
rect 375 2444 395 2496
rect 447 2444 467 2496
rect 519 2444 539 2496
rect 591 2444 611 2496
rect 663 2444 683 2496
rect 735 2444 755 2496
rect 807 2444 827 2496
rect 879 2444 899 2496
rect 951 2444 971 2496
rect 1023 2444 1043 2496
rect 1095 2444 1115 2496
rect 1167 2444 1187 2496
rect 1239 2444 1259 2496
rect 1311 2444 1331 2496
rect 1383 2444 1403 2496
rect 1455 2444 1475 2496
rect 1527 2444 1547 2496
rect 1599 2444 1619 2496
rect 1671 2444 1691 2496
rect 1743 2444 1763 2496
rect 1815 2444 1835 2496
rect 1887 2444 1907 2496
rect 1959 2444 1979 2496
rect 2031 2444 2051 2496
rect 2103 2444 2123 2496
rect 2175 2444 2195 2496
rect 2247 2444 2267 2496
rect 2319 2444 2339 2496
rect 2391 2444 2411 2496
rect 2463 2444 2483 2496
rect 2535 2444 2555 2496
rect 2607 2444 2627 2496
rect 2679 2444 2699 2496
rect 2751 2444 2771 2496
rect 2823 2444 2843 2496
rect 2895 2444 2915 2496
rect 2967 2444 2987 2496
rect 3039 2444 3059 2496
rect 3111 2444 3131 2496
rect 3183 2444 3203 2496
rect 3255 2444 3275 2496
rect 3327 2444 3347 2496
rect 3399 2444 3419 2496
rect 3471 2444 3491 2496
rect 3543 2444 3563 2496
rect 3615 2444 3635 2496
rect 3687 2444 3707 2496
rect 3759 2444 3779 2496
rect 3831 2444 3851 2496
rect 3903 2444 3923 2496
rect 3975 2444 3995 2496
rect 4047 2444 4067 2496
rect 4119 2444 4139 2496
rect 4191 2444 4211 2496
rect 4263 2444 4283 2496
rect 4335 2444 4355 2496
rect 4407 2444 4427 2496
rect 4479 2444 4499 2496
rect 4551 2444 4571 2496
rect 4623 2444 4643 2496
rect 4695 2444 4715 2496
rect 4767 2444 4787 2496
rect 4839 2444 4859 2496
rect 4911 2444 4931 2496
rect 4983 2444 5003 2496
rect 5055 2444 5075 2496
rect 5127 2444 5147 2496
rect 5199 2444 5219 2496
rect 5271 2444 5291 2496
rect 5343 2444 5363 2496
rect 5415 2444 5435 2496
rect 5487 2444 5507 2496
rect 5559 2444 5579 2496
rect 5631 2444 5651 2496
rect 5703 2444 5723 2496
rect 5775 2444 5795 2496
rect 5847 2444 5867 2496
rect 5919 2444 5939 2496
rect 5991 2444 6011 2496
rect 6063 2444 6083 2496
rect 6135 2444 6155 2496
rect 6207 2444 6227 2496
rect 6279 2444 6299 2496
rect 6351 2444 6371 2496
rect 6423 2444 6443 2496
rect 6495 2444 6515 2496
rect 6567 2444 6587 2496
rect 6639 2444 6659 2496
rect 6711 2444 6731 2496
rect 6783 2444 6803 2496
rect 6855 2444 6875 2496
rect 6927 2444 6947 2496
rect 6999 2444 7019 2496
rect 7071 2444 7091 2496
rect 7143 2444 7163 2496
rect 7215 2444 7235 2496
rect 7287 2444 7307 2496
rect 7359 2444 7379 2496
rect 7431 2444 7451 2496
rect 7503 2444 7523 2496
rect 7575 2444 7595 2496
rect 7647 2444 7667 2496
rect 7719 2444 7739 2496
rect 7791 2444 7811 2496
rect 7863 2444 7883 2496
rect 7935 2444 7955 2496
rect 8007 2444 8027 2496
rect 8079 2444 8099 2496
rect 8151 2444 8157 2496
rect 173 2424 8157 2444
rect 173 2372 179 2424
rect 231 2372 251 2424
rect 303 2372 323 2424
rect 375 2372 395 2424
rect 447 2372 467 2424
rect 519 2372 539 2424
rect 591 2372 611 2424
rect 663 2372 683 2424
rect 735 2372 755 2424
rect 807 2372 827 2424
rect 879 2372 899 2424
rect 951 2372 971 2424
rect 1023 2372 1043 2424
rect 1095 2372 1115 2424
rect 1167 2372 1187 2424
rect 1239 2372 1259 2424
rect 1311 2372 1331 2424
rect 1383 2372 1403 2424
rect 1455 2372 1475 2424
rect 1527 2372 1547 2424
rect 1599 2372 1619 2424
rect 1671 2372 1691 2424
rect 1743 2372 1763 2424
rect 1815 2372 1835 2424
rect 1887 2372 1907 2424
rect 1959 2372 1979 2424
rect 2031 2372 2051 2424
rect 2103 2372 2123 2424
rect 2175 2372 2195 2424
rect 2247 2372 2267 2424
rect 2319 2372 2339 2424
rect 2391 2372 2411 2424
rect 2463 2372 2483 2424
rect 2535 2372 2555 2424
rect 2607 2372 2627 2424
rect 2679 2372 2699 2424
rect 2751 2372 2771 2424
rect 2823 2372 2843 2424
rect 2895 2372 2915 2424
rect 2967 2372 2987 2424
rect 3039 2372 3059 2424
rect 3111 2372 3131 2424
rect 3183 2372 3203 2424
rect 3255 2372 3275 2424
rect 3327 2372 3347 2424
rect 3399 2372 3419 2424
rect 3471 2372 3491 2424
rect 3543 2372 3563 2424
rect 3615 2372 3635 2424
rect 3687 2372 3707 2424
rect 3759 2372 3779 2424
rect 3831 2372 3851 2424
rect 3903 2372 3923 2424
rect 3975 2372 3995 2424
rect 4047 2372 4067 2424
rect 4119 2372 4139 2424
rect 4191 2372 4211 2424
rect 4263 2372 4283 2424
rect 4335 2372 4355 2424
rect 4407 2372 4427 2424
rect 4479 2372 4499 2424
rect 4551 2372 4571 2424
rect 4623 2372 4643 2424
rect 4695 2372 4715 2424
rect 4767 2372 4787 2424
rect 4839 2372 4859 2424
rect 4911 2372 4931 2424
rect 4983 2372 5003 2424
rect 5055 2372 5075 2424
rect 5127 2372 5147 2424
rect 5199 2372 5219 2424
rect 5271 2372 5291 2424
rect 5343 2372 5363 2424
rect 5415 2372 5435 2424
rect 5487 2372 5507 2424
rect 5559 2372 5579 2424
rect 5631 2372 5651 2424
rect 5703 2372 5723 2424
rect 5775 2372 5795 2424
rect 5847 2372 5867 2424
rect 5919 2372 5939 2424
rect 5991 2372 6011 2424
rect 6063 2372 6083 2424
rect 6135 2372 6155 2424
rect 6207 2372 6227 2424
rect 6279 2372 6299 2424
rect 6351 2372 6371 2424
rect 6423 2372 6443 2424
rect 6495 2372 6515 2424
rect 6567 2372 6587 2424
rect 6639 2372 6659 2424
rect 6711 2372 6731 2424
rect 6783 2372 6803 2424
rect 6855 2372 6875 2424
rect 6927 2372 6947 2424
rect 6999 2372 7019 2424
rect 7071 2372 7091 2424
rect 7143 2372 7163 2424
rect 7215 2372 7235 2424
rect 7287 2372 7307 2424
rect 7359 2372 7379 2424
rect 7431 2372 7451 2424
rect 7503 2372 7523 2424
rect 7575 2372 7595 2424
rect 7647 2372 7667 2424
rect 7719 2372 7739 2424
rect 7791 2372 7811 2424
rect 7863 2372 7883 2424
rect 7935 2372 7955 2424
rect 8007 2372 8027 2424
rect 8079 2372 8099 2424
rect 8151 2372 8157 2424
rect 173 2352 8157 2372
rect 173 2300 179 2352
rect 231 2300 251 2352
rect 303 2300 323 2352
rect 375 2300 395 2352
rect 447 2300 467 2352
rect 519 2300 539 2352
rect 591 2300 611 2352
rect 663 2300 683 2352
rect 735 2300 755 2352
rect 807 2300 827 2352
rect 879 2300 899 2352
rect 951 2300 971 2352
rect 1023 2300 1043 2352
rect 1095 2300 1115 2352
rect 1167 2300 1187 2352
rect 1239 2300 1259 2352
rect 1311 2300 1331 2352
rect 1383 2300 1403 2352
rect 1455 2300 1475 2352
rect 1527 2300 1547 2352
rect 1599 2300 1619 2352
rect 1671 2300 1691 2352
rect 1743 2300 1763 2352
rect 1815 2300 1835 2352
rect 1887 2300 1907 2352
rect 1959 2300 1979 2352
rect 2031 2300 2051 2352
rect 2103 2300 2123 2352
rect 2175 2300 2195 2352
rect 2247 2300 2267 2352
rect 2319 2300 2339 2352
rect 2391 2300 2411 2352
rect 2463 2300 2483 2352
rect 2535 2300 2555 2352
rect 2607 2300 2627 2352
rect 2679 2300 2699 2352
rect 2751 2300 2771 2352
rect 2823 2300 2843 2352
rect 2895 2300 2915 2352
rect 2967 2300 2987 2352
rect 3039 2300 3059 2352
rect 3111 2300 3131 2352
rect 3183 2300 3203 2352
rect 3255 2300 3275 2352
rect 3327 2300 3347 2352
rect 3399 2300 3419 2352
rect 3471 2300 3491 2352
rect 3543 2300 3563 2352
rect 3615 2300 3635 2352
rect 3687 2300 3707 2352
rect 3759 2300 3779 2352
rect 3831 2300 3851 2352
rect 3903 2300 3923 2352
rect 3975 2300 3995 2352
rect 4047 2300 4067 2352
rect 4119 2300 4139 2352
rect 4191 2300 4211 2352
rect 4263 2300 4283 2352
rect 4335 2300 4355 2352
rect 4407 2300 4427 2352
rect 4479 2300 4499 2352
rect 4551 2300 4571 2352
rect 4623 2300 4643 2352
rect 4695 2300 4715 2352
rect 4767 2300 4787 2352
rect 4839 2300 4859 2352
rect 4911 2300 4931 2352
rect 4983 2300 5003 2352
rect 5055 2300 5075 2352
rect 5127 2300 5147 2352
rect 5199 2300 5219 2352
rect 5271 2300 5291 2352
rect 5343 2300 5363 2352
rect 5415 2300 5435 2352
rect 5487 2300 5507 2352
rect 5559 2300 5579 2352
rect 5631 2300 5651 2352
rect 5703 2300 5723 2352
rect 5775 2300 5795 2352
rect 5847 2300 5867 2352
rect 5919 2300 5939 2352
rect 5991 2300 6011 2352
rect 6063 2300 6083 2352
rect 6135 2300 6155 2352
rect 6207 2300 6227 2352
rect 6279 2300 6299 2352
rect 6351 2300 6371 2352
rect 6423 2300 6443 2352
rect 6495 2300 6515 2352
rect 6567 2300 6587 2352
rect 6639 2300 6659 2352
rect 6711 2300 6731 2352
rect 6783 2300 6803 2352
rect 6855 2300 6875 2352
rect 6927 2300 6947 2352
rect 6999 2300 7019 2352
rect 7071 2300 7091 2352
rect 7143 2300 7163 2352
rect 7215 2300 7235 2352
rect 7287 2300 7307 2352
rect 7359 2300 7379 2352
rect 7431 2300 7451 2352
rect 7503 2300 7523 2352
rect 7575 2300 7595 2352
rect 7647 2300 7667 2352
rect 7719 2300 7739 2352
rect 7791 2300 7811 2352
rect 7863 2300 7883 2352
rect 7935 2300 7955 2352
rect 8007 2300 8027 2352
rect 8079 2300 8099 2352
rect 8151 2300 8157 2352
rect 173 2294 8157 2300
rect 180 162 318 168
rect 180 110 186 162
rect 238 110 260 162
rect 312 110 318 162
rect 180 88 318 110
rect 180 36 186 88
rect 238 36 260 88
rect 312 36 318 88
rect 180 30 318 36
use nfet$1  nfet$1_0
timestamp 1698982078
transform 0 -1 6205 1 0 282
box -1 0 715 6146
use nfet$2  nfet$2_0
timestamp 1698982078
transform 0 -1 389 -1 0 300
box -1 0 301 346
use pfet  pfet_0
timestamp 1698982078
transform 0 -1 8241 1 0 996
box 0 0 1595 8220
<< labels >>
flabel metal1 s 18 137 134 250 0 FreeSans 44 0 0 0 CTRL
port 2 nsew
flabel metal1 s 176 846 8154 1254 0 FreeSans 44 0 0 0 OUT
port 3 nsew
flabel metal1 s 266 1067 266 1067 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 4296 1065 4296 1065 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 6363 1072 6363 1072 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 2054 1101 2054 1101 0 FreeSans 44 0 0 0 OUT
flabel metal1 s 0 466 115 2050 0 FreeSans 44 0 0 0 IN
port 4 nsew
flabel metal1 s 55 491 55 491 0 FreeSans 44 0 0 0 IN
flabel metal1 s 56 1378 56 1378 0 FreeSans 44 0 0 0 IN
flabel metal1 s 56 1745 56 1745 0 FreeSans 44 0 0 0 IN
flabel metal1 s 58 992 58 992 0 FreeSans 44 0 0 0 IN
flabel metal2 s 180 30 318 168 0 FreeSans 44 0 0 0 VSS
port 6 nsew
flabel metal2 s 173 2294 8157 2502 0 FreeSans 44 0 0 0 VDD
port 7 nsew
flabel metal2 s 8112 2401 8112 2401 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 4127 2395 4127 2395 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 6470 2387 6470 2387 0 FreeSans 44 0 0 0 VDD
flabel metal2 s 2102 2408 2102 2408 0 FreeSans 44 0 0 0 VDD
<< end >>
