magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -350 -90 7270 25260
<< l68d20 >>
rect 3970 2796 6760 4979
rect 2700 5281 6760 7464
rect 1430 7766 6760 9949
rect 160 10251 6760 12434
rect 160 12736 6760 14919
rect 1430 15221 6760 17404
rect 2700 17706 6760 19889
rect 3970 20191 6760 22374
rect 160 15471 410 17575
rect 5205 135 5525 2255
rect 5205 22670 5525 24790
<< l68d16 >>
rect 3970 140 4220 2244
rect 2700 2625 2950 4729
rect 1430 5110 1680 7214
rect 160 7595 410 9699
rect 160 15471 410 17575
rect 1430 17956 1680 20060
rect 2700 20441 2950 22545
rect 3970 22926 4220 25030
rect 3970 20191 6760 22374
<< l68d44 >>
rect 5290 1660 5440 1810
rect 5290 1300 5440 1450
rect 5290 940 5440 1090
rect 5290 580 5440 730
rect 5290 220 5440 370
rect 5290 24195 5440 24345
rect 5290 23835 5440 23985
rect 5290 23475 5440 23625
rect 5290 23115 5440 23265
rect 5290 22755 5440 22905
rect 5290 2021 5440 2171
rect 5290 24555 5440 24705
<< l69d20 >>
rect 5205 135 5525 2256
rect 5205 22670 5525 24790
<< l69d16 >>
rect 5205 135 5525 2256
rect 5205 22670 5525 24790
<< labels >>
rlabel l68d5 4667 20363 4667 20363 0 OUT
rlabel l68d5 4686 21303 4686 21303 0 OUT
rlabel l68d5 4617 22248 4617 22248 0 OUT
rlabel l68d5 1543 18113 1543 18113 0 DAC5
rlabel l68d5 1556 19023 1556 19023 0 DAC5
rlabel l68d5 1543 19921 1543 19921 0 DAC5
rlabel l68d5 2823 20590 2823 20590 0 DAC6
rlabel l68d5 4088 24886 4088 24886 0 DAC7
rlabel l68d5 2815 22406 2815 22406 0 DAC6
rlabel l68d5 2827 21484 2827 21484 0 DAC6
rlabel l68d5 4088 23079 4088 23079 0 DAC7
rlabel l68d5 4085 23984 4085 23984 0 DAC7
rlabel l68d5 5984 22193 5984 22193 0 OUT
rlabel l68d5 5979 21367 5979 21367 0 OUT
rlabel l68d5 5984 20400 5984 20400 0 OUT
rlabel l68d5 284 17415 284 17415 0 DAC4
rlabel l68d5 276 16522 276 16522 0 DAC4
rlabel l68d5 276 15624 276 15624 0 DAC4
rlabel l68d5 288 9569 288 9569 0 DAC3
rlabel l68d5 293 8679 293 8679 0 DAC3
rlabel l68d5 280 7753 280 7753 0 DAC3
rlabel l68d5 1561 6190 1561 6190 0 DAC2
rlabel l68d5 1547 7056 1547 7056 0 DAC2
rlabel l68d5 1561 5274 1561 5274 0 DAC2
rlabel l68d5 2824 3692 2824 3692 0 DAC1
rlabel l68d5 2841 4597 2841 4597 0 DAC1
rlabel l68d5 2830 2782 2830 2782 0 DAC1
rlabel l68d5 4107 1204 4107 1204 0 DAC0
rlabel l68d5 4092 2096 4092 2096 0 DAC0
rlabel l68d5 4092 298 4092 298 0 DAC0
rlabel l69d5 5360 24650 5360 24650 0 VDD
rlabel l69d5 5360 23746 5360 23746 0 VDD
rlabel l69d5 5360 22827 5360 22827 0 VDD
rlabel l69d5 5369 1194 5369 1194 0 VSS
rlabel l69d5 5351 289 5351 289 0 VSS
rlabel l69d5 5359 2092 5359 2092 0 VSS
use res_polyx243 res_polyx243_1
timestamp 1698899266
transform 1 0 285 0 1 15195
box -635 -2610 635 2610
use res_polyx243 res_polyx243_2
timestamp 1698899266
transform 1 0 1555 0 1 7490
box -635 -2610 635 2610
use res_polyx244 res_polyx244_1
timestamp 1698899266
transform 1 0 5365 0 1 12585
box -635 -2485 635 2485
use res_polyx243 res_polyx243_3
timestamp 1698899266
transform 1 0 1555 0 1 17680
box -635 -2610 635 2610
use res_polyx243 res_polyx243_4
timestamp 1698899266
transform 1 0 285 0 1 9975
box -635 -2610 635 2610
use res_polyx243 res_polyx243_5
timestamp 1698899266
transform 1 0 5365 0 1 2520
box -635 -2610 635 2610
use res_polyx244 res_polyx244_2
timestamp 1698899266
transform 1 0 5365 0 1 7615
box -635 -2485 635 2485
use res_polyx244 res_polyx244_3
timestamp 1698899266
transform 1 0 6635 0 1 5130
box -635 -2485 635 2485
use res_polyx244 res_polyx244_4
timestamp 1698899266
transform 1 0 6635 0 1 15070
box -635 -2485 635 2485
use res_polyx243 res_polyx243_6
timestamp 1698899266
transform 1 0 4095 0 1 22650
box -635 -2610 635 2610
use res_polyx244 res_polyx244_5
timestamp 1698899266
transform 1 0 6635 0 1 20040
box -635 -2485 635 2485
use res_polyx243 res_polyx243_7
timestamp 1698899266
transform 1 0 2825 0 1 20165
box -635 -2610 635 2610
use res_polyx244 res_polyx244_6
timestamp 1698899266
transform 1 0 5365 0 1 17555
box -635 -2485 635 2485
use res_polyx244 res_polyx244_7
timestamp 1698899266
transform 1 0 5365 0 1 22525
box -635 -2485 635 2485
use res_polyx243 res_polyx243_8
timestamp 1698899266
transform 1 0 4095 0 1 2520
box -635 -2610 635 2610
use res_polyx243 res_polyx243_9
timestamp 1698899266
transform 1 0 2825 0 1 5005
box -635 -2610 635 2610
use res_polyx244 res_polyx244_8
timestamp 1698899266
transform 1 0 6635 0 1 10100
box -635 -2485 635 2485
<< end >>
