magic
tech sky130A
magscale 1 2
timestamp 1699066547
<< pwell >>
rect -1 14 715 6066
<< nmos >>
rect 157 40 557 6040
<< ndiff >>
rect 25 6009 157 6040
rect 25 5975 38 6009
rect 72 5975 110 6009
rect 144 5975 157 6009
rect 25 5937 157 5975
rect 25 5903 38 5937
rect 72 5903 110 5937
rect 144 5903 157 5937
rect 25 5865 157 5903
rect 25 5831 38 5865
rect 72 5831 110 5865
rect 144 5831 157 5865
rect 25 5793 157 5831
rect 25 5759 38 5793
rect 72 5759 110 5793
rect 144 5759 157 5793
rect 25 5721 157 5759
rect 25 5687 38 5721
rect 72 5687 110 5721
rect 144 5687 157 5721
rect 25 5649 157 5687
rect 25 5615 38 5649
rect 72 5615 110 5649
rect 144 5615 157 5649
rect 25 5577 157 5615
rect 25 5543 38 5577
rect 72 5543 110 5577
rect 144 5543 157 5577
rect 25 5505 157 5543
rect 25 5471 38 5505
rect 72 5471 110 5505
rect 144 5471 157 5505
rect 25 5433 157 5471
rect 25 5399 38 5433
rect 72 5399 110 5433
rect 144 5399 157 5433
rect 25 5361 157 5399
rect 25 5327 38 5361
rect 72 5327 110 5361
rect 144 5327 157 5361
rect 25 5289 157 5327
rect 25 5255 38 5289
rect 72 5255 110 5289
rect 144 5255 157 5289
rect 25 5217 157 5255
rect 25 5183 38 5217
rect 72 5183 110 5217
rect 144 5183 157 5217
rect 25 5145 157 5183
rect 25 5111 38 5145
rect 72 5111 110 5145
rect 144 5111 157 5145
rect 25 5073 157 5111
rect 25 5039 38 5073
rect 72 5039 110 5073
rect 144 5039 157 5073
rect 25 5001 157 5039
rect 25 4967 38 5001
rect 72 4967 110 5001
rect 144 4967 157 5001
rect 25 4929 157 4967
rect 25 4895 38 4929
rect 72 4895 110 4929
rect 144 4895 157 4929
rect 25 4857 157 4895
rect 25 4823 38 4857
rect 72 4823 110 4857
rect 144 4823 157 4857
rect 25 4785 157 4823
rect 25 4751 38 4785
rect 72 4751 110 4785
rect 144 4751 157 4785
rect 25 4713 157 4751
rect 25 4679 38 4713
rect 72 4679 110 4713
rect 144 4679 157 4713
rect 25 4641 157 4679
rect 25 4607 38 4641
rect 72 4607 110 4641
rect 144 4607 157 4641
rect 25 4569 157 4607
rect 25 4535 38 4569
rect 72 4535 110 4569
rect 144 4535 157 4569
rect 25 4497 157 4535
rect 25 4463 38 4497
rect 72 4463 110 4497
rect 144 4463 157 4497
rect 25 4425 157 4463
rect 25 4391 38 4425
rect 72 4391 110 4425
rect 144 4391 157 4425
rect 25 4353 157 4391
rect 25 4319 38 4353
rect 72 4319 110 4353
rect 144 4319 157 4353
rect 25 4281 157 4319
rect 25 4247 38 4281
rect 72 4247 110 4281
rect 144 4247 157 4281
rect 25 4209 157 4247
rect 25 4175 38 4209
rect 72 4175 110 4209
rect 144 4175 157 4209
rect 25 4137 157 4175
rect 25 4103 38 4137
rect 72 4103 110 4137
rect 144 4103 157 4137
rect 25 4065 157 4103
rect 25 4031 38 4065
rect 72 4031 110 4065
rect 144 4031 157 4065
rect 25 3993 157 4031
rect 25 3959 38 3993
rect 72 3959 110 3993
rect 144 3959 157 3993
rect 25 3921 157 3959
rect 25 3887 38 3921
rect 72 3887 110 3921
rect 144 3887 157 3921
rect 25 3849 157 3887
rect 25 3815 38 3849
rect 72 3815 110 3849
rect 144 3815 157 3849
rect 25 3777 157 3815
rect 25 3743 38 3777
rect 72 3743 110 3777
rect 144 3743 157 3777
rect 25 3705 157 3743
rect 25 3671 38 3705
rect 72 3671 110 3705
rect 144 3671 157 3705
rect 25 3633 157 3671
rect 25 3599 38 3633
rect 72 3599 110 3633
rect 144 3599 157 3633
rect 25 3561 157 3599
rect 25 3527 38 3561
rect 72 3527 110 3561
rect 144 3527 157 3561
rect 25 3489 157 3527
rect 25 3455 38 3489
rect 72 3455 110 3489
rect 144 3455 157 3489
rect 25 3417 157 3455
rect 25 3383 38 3417
rect 72 3383 110 3417
rect 144 3383 157 3417
rect 25 3345 157 3383
rect 25 3311 38 3345
rect 72 3311 110 3345
rect 144 3311 157 3345
rect 25 3273 157 3311
rect 25 3239 38 3273
rect 72 3239 110 3273
rect 144 3239 157 3273
rect 25 3201 157 3239
rect 25 3167 38 3201
rect 72 3167 110 3201
rect 144 3167 157 3201
rect 25 3129 157 3167
rect 25 3095 38 3129
rect 72 3095 110 3129
rect 144 3095 157 3129
rect 25 3057 157 3095
rect 25 3023 38 3057
rect 72 3023 110 3057
rect 144 3023 157 3057
rect 25 2985 157 3023
rect 25 2951 38 2985
rect 72 2951 110 2985
rect 144 2951 157 2985
rect 25 2913 157 2951
rect 25 2879 38 2913
rect 72 2879 110 2913
rect 144 2879 157 2913
rect 25 2841 157 2879
rect 25 2807 38 2841
rect 72 2807 110 2841
rect 144 2807 157 2841
rect 25 2769 157 2807
rect 25 2735 38 2769
rect 72 2735 110 2769
rect 144 2735 157 2769
rect 25 2697 157 2735
rect 25 2663 38 2697
rect 72 2663 110 2697
rect 144 2663 157 2697
rect 25 2625 157 2663
rect 25 2591 38 2625
rect 72 2591 110 2625
rect 144 2591 157 2625
rect 25 2553 157 2591
rect 25 2519 38 2553
rect 72 2519 110 2553
rect 144 2519 157 2553
rect 25 2481 157 2519
rect 25 2447 38 2481
rect 72 2447 110 2481
rect 144 2447 157 2481
rect 25 2409 157 2447
rect 25 2375 38 2409
rect 72 2375 110 2409
rect 144 2375 157 2409
rect 25 2337 157 2375
rect 25 2303 38 2337
rect 72 2303 110 2337
rect 144 2303 157 2337
rect 25 2265 157 2303
rect 25 2231 38 2265
rect 72 2231 110 2265
rect 144 2231 157 2265
rect 25 2193 157 2231
rect 25 2159 38 2193
rect 72 2159 110 2193
rect 144 2159 157 2193
rect 25 2121 157 2159
rect 25 2087 38 2121
rect 72 2087 110 2121
rect 144 2087 157 2121
rect 25 2049 157 2087
rect 25 2015 38 2049
rect 72 2015 110 2049
rect 144 2015 157 2049
rect 25 1977 157 2015
rect 25 1943 38 1977
rect 72 1943 110 1977
rect 144 1943 157 1977
rect 25 1905 157 1943
rect 25 1871 38 1905
rect 72 1871 110 1905
rect 144 1871 157 1905
rect 25 1833 157 1871
rect 25 1799 38 1833
rect 72 1799 110 1833
rect 144 1799 157 1833
rect 25 1761 157 1799
rect 25 1727 38 1761
rect 72 1727 110 1761
rect 144 1727 157 1761
rect 25 1689 157 1727
rect 25 1655 38 1689
rect 72 1655 110 1689
rect 144 1655 157 1689
rect 25 1617 157 1655
rect 25 1583 38 1617
rect 72 1583 110 1617
rect 144 1583 157 1617
rect 25 1545 157 1583
rect 25 1511 38 1545
rect 72 1511 110 1545
rect 144 1511 157 1545
rect 25 1473 157 1511
rect 25 1439 38 1473
rect 72 1439 110 1473
rect 144 1439 157 1473
rect 25 1401 157 1439
rect 25 1367 38 1401
rect 72 1367 110 1401
rect 144 1367 157 1401
rect 25 1329 157 1367
rect 25 1295 38 1329
rect 72 1295 110 1329
rect 144 1295 157 1329
rect 25 1257 157 1295
rect 25 1223 38 1257
rect 72 1223 110 1257
rect 144 1223 157 1257
rect 25 1185 157 1223
rect 25 1151 38 1185
rect 72 1151 110 1185
rect 144 1151 157 1185
rect 25 1113 157 1151
rect 25 1079 38 1113
rect 72 1079 110 1113
rect 144 1079 157 1113
rect 25 1041 157 1079
rect 25 1007 38 1041
rect 72 1007 110 1041
rect 144 1007 157 1041
rect 25 969 157 1007
rect 25 935 38 969
rect 72 935 110 969
rect 144 935 157 969
rect 25 897 157 935
rect 25 863 38 897
rect 72 863 110 897
rect 144 863 157 897
rect 25 825 157 863
rect 25 791 38 825
rect 72 791 110 825
rect 144 791 157 825
rect 25 753 157 791
rect 25 719 38 753
rect 72 719 110 753
rect 144 719 157 753
rect 25 681 157 719
rect 25 647 38 681
rect 72 647 110 681
rect 144 647 157 681
rect 25 609 157 647
rect 25 575 38 609
rect 72 575 110 609
rect 144 575 157 609
rect 25 537 157 575
rect 25 503 38 537
rect 72 503 110 537
rect 144 503 157 537
rect 25 465 157 503
rect 25 431 38 465
rect 72 431 110 465
rect 144 431 157 465
rect 25 393 157 431
rect 25 359 38 393
rect 72 359 110 393
rect 144 359 157 393
rect 25 321 157 359
rect 25 287 38 321
rect 72 287 110 321
rect 144 287 157 321
rect 25 249 157 287
rect 25 215 38 249
rect 72 215 110 249
rect 144 215 157 249
rect 25 177 157 215
rect 25 143 38 177
rect 72 143 110 177
rect 144 143 157 177
rect 25 105 157 143
rect 25 71 38 105
rect 72 71 110 105
rect 144 71 157 105
rect 25 40 157 71
rect 557 6009 689 6040
rect 557 5975 570 6009
rect 604 5975 642 6009
rect 676 5975 689 6009
rect 557 5937 689 5975
rect 557 5903 570 5937
rect 604 5903 642 5937
rect 676 5903 689 5937
rect 557 5865 689 5903
rect 557 5831 570 5865
rect 604 5831 642 5865
rect 676 5831 689 5865
rect 557 5793 689 5831
rect 557 5759 570 5793
rect 604 5759 642 5793
rect 676 5759 689 5793
rect 557 5721 689 5759
rect 557 5687 570 5721
rect 604 5687 642 5721
rect 676 5687 689 5721
rect 557 5649 689 5687
rect 557 5615 570 5649
rect 604 5615 642 5649
rect 676 5615 689 5649
rect 557 5577 689 5615
rect 557 5543 570 5577
rect 604 5543 642 5577
rect 676 5543 689 5577
rect 557 5505 689 5543
rect 557 5471 570 5505
rect 604 5471 642 5505
rect 676 5471 689 5505
rect 557 5433 689 5471
rect 557 5399 570 5433
rect 604 5399 642 5433
rect 676 5399 689 5433
rect 557 5361 689 5399
rect 557 5327 570 5361
rect 604 5327 642 5361
rect 676 5327 689 5361
rect 557 5289 689 5327
rect 557 5255 570 5289
rect 604 5255 642 5289
rect 676 5255 689 5289
rect 557 5217 689 5255
rect 557 5183 570 5217
rect 604 5183 642 5217
rect 676 5183 689 5217
rect 557 5145 689 5183
rect 557 5111 570 5145
rect 604 5111 642 5145
rect 676 5111 689 5145
rect 557 5073 689 5111
rect 557 5039 570 5073
rect 604 5039 642 5073
rect 676 5039 689 5073
rect 557 5001 689 5039
rect 557 4967 570 5001
rect 604 4967 642 5001
rect 676 4967 689 5001
rect 557 4929 689 4967
rect 557 4895 570 4929
rect 604 4895 642 4929
rect 676 4895 689 4929
rect 557 4857 689 4895
rect 557 4823 570 4857
rect 604 4823 642 4857
rect 676 4823 689 4857
rect 557 4785 689 4823
rect 557 4751 570 4785
rect 604 4751 642 4785
rect 676 4751 689 4785
rect 557 4713 689 4751
rect 557 4679 570 4713
rect 604 4679 642 4713
rect 676 4679 689 4713
rect 557 4641 689 4679
rect 557 4607 570 4641
rect 604 4607 642 4641
rect 676 4607 689 4641
rect 557 4569 689 4607
rect 557 4535 570 4569
rect 604 4535 642 4569
rect 676 4535 689 4569
rect 557 4497 689 4535
rect 557 4463 570 4497
rect 604 4463 642 4497
rect 676 4463 689 4497
rect 557 4425 689 4463
rect 557 4391 570 4425
rect 604 4391 642 4425
rect 676 4391 689 4425
rect 557 4353 689 4391
rect 557 4319 570 4353
rect 604 4319 642 4353
rect 676 4319 689 4353
rect 557 4281 689 4319
rect 557 4247 570 4281
rect 604 4247 642 4281
rect 676 4247 689 4281
rect 557 4209 689 4247
rect 557 4175 570 4209
rect 604 4175 642 4209
rect 676 4175 689 4209
rect 557 4137 689 4175
rect 557 4103 570 4137
rect 604 4103 642 4137
rect 676 4103 689 4137
rect 557 4065 689 4103
rect 557 4031 570 4065
rect 604 4031 642 4065
rect 676 4031 689 4065
rect 557 3993 689 4031
rect 557 3959 570 3993
rect 604 3959 642 3993
rect 676 3959 689 3993
rect 557 3921 689 3959
rect 557 3887 570 3921
rect 604 3887 642 3921
rect 676 3887 689 3921
rect 557 3849 689 3887
rect 557 3815 570 3849
rect 604 3815 642 3849
rect 676 3815 689 3849
rect 557 3777 689 3815
rect 557 3743 570 3777
rect 604 3743 642 3777
rect 676 3743 689 3777
rect 557 3705 689 3743
rect 557 3671 570 3705
rect 604 3671 642 3705
rect 676 3671 689 3705
rect 557 3633 689 3671
rect 557 3599 570 3633
rect 604 3599 642 3633
rect 676 3599 689 3633
rect 557 3561 689 3599
rect 557 3527 570 3561
rect 604 3527 642 3561
rect 676 3527 689 3561
rect 557 3489 689 3527
rect 557 3455 570 3489
rect 604 3455 642 3489
rect 676 3455 689 3489
rect 557 3417 689 3455
rect 557 3383 570 3417
rect 604 3383 642 3417
rect 676 3383 689 3417
rect 557 3345 689 3383
rect 557 3311 570 3345
rect 604 3311 642 3345
rect 676 3311 689 3345
rect 557 3273 689 3311
rect 557 3239 570 3273
rect 604 3239 642 3273
rect 676 3239 689 3273
rect 557 3201 689 3239
rect 557 3167 570 3201
rect 604 3167 642 3201
rect 676 3167 689 3201
rect 557 3129 689 3167
rect 557 3095 570 3129
rect 604 3095 642 3129
rect 676 3095 689 3129
rect 557 3057 689 3095
rect 557 3023 570 3057
rect 604 3023 642 3057
rect 676 3023 689 3057
rect 557 2985 689 3023
rect 557 2951 570 2985
rect 604 2951 642 2985
rect 676 2951 689 2985
rect 557 2913 689 2951
rect 557 2879 570 2913
rect 604 2879 642 2913
rect 676 2879 689 2913
rect 557 2841 689 2879
rect 557 2807 570 2841
rect 604 2807 642 2841
rect 676 2807 689 2841
rect 557 2769 689 2807
rect 557 2735 570 2769
rect 604 2735 642 2769
rect 676 2735 689 2769
rect 557 2697 689 2735
rect 557 2663 570 2697
rect 604 2663 642 2697
rect 676 2663 689 2697
rect 557 2625 689 2663
rect 557 2591 570 2625
rect 604 2591 642 2625
rect 676 2591 689 2625
rect 557 2553 689 2591
rect 557 2519 570 2553
rect 604 2519 642 2553
rect 676 2519 689 2553
rect 557 2481 689 2519
rect 557 2447 570 2481
rect 604 2447 642 2481
rect 676 2447 689 2481
rect 557 2409 689 2447
rect 557 2375 570 2409
rect 604 2375 642 2409
rect 676 2375 689 2409
rect 557 2337 689 2375
rect 557 2303 570 2337
rect 604 2303 642 2337
rect 676 2303 689 2337
rect 557 2265 689 2303
rect 557 2231 570 2265
rect 604 2231 642 2265
rect 676 2231 689 2265
rect 557 2193 689 2231
rect 557 2159 570 2193
rect 604 2159 642 2193
rect 676 2159 689 2193
rect 557 2121 689 2159
rect 557 2087 570 2121
rect 604 2087 642 2121
rect 676 2087 689 2121
rect 557 2049 689 2087
rect 557 2015 570 2049
rect 604 2015 642 2049
rect 676 2015 689 2049
rect 557 1977 689 2015
rect 557 1943 570 1977
rect 604 1943 642 1977
rect 676 1943 689 1977
rect 557 1905 689 1943
rect 557 1871 570 1905
rect 604 1871 642 1905
rect 676 1871 689 1905
rect 557 1833 689 1871
rect 557 1799 570 1833
rect 604 1799 642 1833
rect 676 1799 689 1833
rect 557 1761 689 1799
rect 557 1727 570 1761
rect 604 1727 642 1761
rect 676 1727 689 1761
rect 557 1689 689 1727
rect 557 1655 570 1689
rect 604 1655 642 1689
rect 676 1655 689 1689
rect 557 1617 689 1655
rect 557 1583 570 1617
rect 604 1583 642 1617
rect 676 1583 689 1617
rect 557 1545 689 1583
rect 557 1511 570 1545
rect 604 1511 642 1545
rect 676 1511 689 1545
rect 557 1473 689 1511
rect 557 1439 570 1473
rect 604 1439 642 1473
rect 676 1439 689 1473
rect 557 1401 689 1439
rect 557 1367 570 1401
rect 604 1367 642 1401
rect 676 1367 689 1401
rect 557 1329 689 1367
rect 557 1295 570 1329
rect 604 1295 642 1329
rect 676 1295 689 1329
rect 557 1257 689 1295
rect 557 1223 570 1257
rect 604 1223 642 1257
rect 676 1223 689 1257
rect 557 1185 689 1223
rect 557 1151 570 1185
rect 604 1151 642 1185
rect 676 1151 689 1185
rect 557 1113 689 1151
rect 557 1079 570 1113
rect 604 1079 642 1113
rect 676 1079 689 1113
rect 557 1041 689 1079
rect 557 1007 570 1041
rect 604 1007 642 1041
rect 676 1007 689 1041
rect 557 969 689 1007
rect 557 935 570 969
rect 604 935 642 969
rect 676 935 689 969
rect 557 897 689 935
rect 557 863 570 897
rect 604 863 642 897
rect 676 863 689 897
rect 557 825 689 863
rect 557 791 570 825
rect 604 791 642 825
rect 676 791 689 825
rect 557 753 689 791
rect 557 719 570 753
rect 604 719 642 753
rect 676 719 689 753
rect 557 681 689 719
rect 557 647 570 681
rect 604 647 642 681
rect 676 647 689 681
rect 557 609 689 647
rect 557 575 570 609
rect 604 575 642 609
rect 676 575 689 609
rect 557 537 689 575
rect 557 503 570 537
rect 604 503 642 537
rect 676 503 689 537
rect 557 465 689 503
rect 557 431 570 465
rect 604 431 642 465
rect 676 431 689 465
rect 557 393 689 431
rect 557 359 570 393
rect 604 359 642 393
rect 676 359 689 393
rect 557 321 689 359
rect 557 287 570 321
rect 604 287 642 321
rect 676 287 689 321
rect 557 249 689 287
rect 557 215 570 249
rect 604 215 642 249
rect 676 215 689 249
rect 557 177 689 215
rect 557 143 570 177
rect 604 143 642 177
rect 676 143 689 177
rect 557 105 689 143
rect 557 71 570 105
rect 604 71 642 105
rect 676 71 689 105
rect 557 40 689 71
<< ndiffc >>
rect 38 5975 72 6009
rect 110 5975 144 6009
rect 38 5903 72 5937
rect 110 5903 144 5937
rect 38 5831 72 5865
rect 110 5831 144 5865
rect 38 5759 72 5793
rect 110 5759 144 5793
rect 38 5687 72 5721
rect 110 5687 144 5721
rect 38 5615 72 5649
rect 110 5615 144 5649
rect 38 5543 72 5577
rect 110 5543 144 5577
rect 38 5471 72 5505
rect 110 5471 144 5505
rect 38 5399 72 5433
rect 110 5399 144 5433
rect 38 5327 72 5361
rect 110 5327 144 5361
rect 38 5255 72 5289
rect 110 5255 144 5289
rect 38 5183 72 5217
rect 110 5183 144 5217
rect 38 5111 72 5145
rect 110 5111 144 5145
rect 38 5039 72 5073
rect 110 5039 144 5073
rect 38 4967 72 5001
rect 110 4967 144 5001
rect 38 4895 72 4929
rect 110 4895 144 4929
rect 38 4823 72 4857
rect 110 4823 144 4857
rect 38 4751 72 4785
rect 110 4751 144 4785
rect 38 4679 72 4713
rect 110 4679 144 4713
rect 38 4607 72 4641
rect 110 4607 144 4641
rect 38 4535 72 4569
rect 110 4535 144 4569
rect 38 4463 72 4497
rect 110 4463 144 4497
rect 38 4391 72 4425
rect 110 4391 144 4425
rect 38 4319 72 4353
rect 110 4319 144 4353
rect 38 4247 72 4281
rect 110 4247 144 4281
rect 38 4175 72 4209
rect 110 4175 144 4209
rect 38 4103 72 4137
rect 110 4103 144 4137
rect 38 4031 72 4065
rect 110 4031 144 4065
rect 38 3959 72 3993
rect 110 3959 144 3993
rect 38 3887 72 3921
rect 110 3887 144 3921
rect 38 3815 72 3849
rect 110 3815 144 3849
rect 38 3743 72 3777
rect 110 3743 144 3777
rect 38 3671 72 3705
rect 110 3671 144 3705
rect 38 3599 72 3633
rect 110 3599 144 3633
rect 38 3527 72 3561
rect 110 3527 144 3561
rect 38 3455 72 3489
rect 110 3455 144 3489
rect 38 3383 72 3417
rect 110 3383 144 3417
rect 38 3311 72 3345
rect 110 3311 144 3345
rect 38 3239 72 3273
rect 110 3239 144 3273
rect 38 3167 72 3201
rect 110 3167 144 3201
rect 38 3095 72 3129
rect 110 3095 144 3129
rect 38 3023 72 3057
rect 110 3023 144 3057
rect 38 2951 72 2985
rect 110 2951 144 2985
rect 38 2879 72 2913
rect 110 2879 144 2913
rect 38 2807 72 2841
rect 110 2807 144 2841
rect 38 2735 72 2769
rect 110 2735 144 2769
rect 38 2663 72 2697
rect 110 2663 144 2697
rect 38 2591 72 2625
rect 110 2591 144 2625
rect 38 2519 72 2553
rect 110 2519 144 2553
rect 38 2447 72 2481
rect 110 2447 144 2481
rect 38 2375 72 2409
rect 110 2375 144 2409
rect 38 2303 72 2337
rect 110 2303 144 2337
rect 38 2231 72 2265
rect 110 2231 144 2265
rect 38 2159 72 2193
rect 110 2159 144 2193
rect 38 2087 72 2121
rect 110 2087 144 2121
rect 38 2015 72 2049
rect 110 2015 144 2049
rect 38 1943 72 1977
rect 110 1943 144 1977
rect 38 1871 72 1905
rect 110 1871 144 1905
rect 38 1799 72 1833
rect 110 1799 144 1833
rect 38 1727 72 1761
rect 110 1727 144 1761
rect 38 1655 72 1689
rect 110 1655 144 1689
rect 38 1583 72 1617
rect 110 1583 144 1617
rect 38 1511 72 1545
rect 110 1511 144 1545
rect 38 1439 72 1473
rect 110 1439 144 1473
rect 38 1367 72 1401
rect 110 1367 144 1401
rect 38 1295 72 1329
rect 110 1295 144 1329
rect 38 1223 72 1257
rect 110 1223 144 1257
rect 38 1151 72 1185
rect 110 1151 144 1185
rect 38 1079 72 1113
rect 110 1079 144 1113
rect 38 1007 72 1041
rect 110 1007 144 1041
rect 38 935 72 969
rect 110 935 144 969
rect 38 863 72 897
rect 110 863 144 897
rect 38 791 72 825
rect 110 791 144 825
rect 38 719 72 753
rect 110 719 144 753
rect 38 647 72 681
rect 110 647 144 681
rect 38 575 72 609
rect 110 575 144 609
rect 38 503 72 537
rect 110 503 144 537
rect 38 431 72 465
rect 110 431 144 465
rect 38 359 72 393
rect 110 359 144 393
rect 38 287 72 321
rect 110 287 144 321
rect 38 215 72 249
rect 110 215 144 249
rect 38 143 72 177
rect 110 143 144 177
rect 38 71 72 105
rect 110 71 144 105
rect 570 5975 604 6009
rect 642 5975 676 6009
rect 570 5903 604 5937
rect 642 5903 676 5937
rect 570 5831 604 5865
rect 642 5831 676 5865
rect 570 5759 604 5793
rect 642 5759 676 5793
rect 570 5687 604 5721
rect 642 5687 676 5721
rect 570 5615 604 5649
rect 642 5615 676 5649
rect 570 5543 604 5577
rect 642 5543 676 5577
rect 570 5471 604 5505
rect 642 5471 676 5505
rect 570 5399 604 5433
rect 642 5399 676 5433
rect 570 5327 604 5361
rect 642 5327 676 5361
rect 570 5255 604 5289
rect 642 5255 676 5289
rect 570 5183 604 5217
rect 642 5183 676 5217
rect 570 5111 604 5145
rect 642 5111 676 5145
rect 570 5039 604 5073
rect 642 5039 676 5073
rect 570 4967 604 5001
rect 642 4967 676 5001
rect 570 4895 604 4929
rect 642 4895 676 4929
rect 570 4823 604 4857
rect 642 4823 676 4857
rect 570 4751 604 4785
rect 642 4751 676 4785
rect 570 4679 604 4713
rect 642 4679 676 4713
rect 570 4607 604 4641
rect 642 4607 676 4641
rect 570 4535 604 4569
rect 642 4535 676 4569
rect 570 4463 604 4497
rect 642 4463 676 4497
rect 570 4391 604 4425
rect 642 4391 676 4425
rect 570 4319 604 4353
rect 642 4319 676 4353
rect 570 4247 604 4281
rect 642 4247 676 4281
rect 570 4175 604 4209
rect 642 4175 676 4209
rect 570 4103 604 4137
rect 642 4103 676 4137
rect 570 4031 604 4065
rect 642 4031 676 4065
rect 570 3959 604 3993
rect 642 3959 676 3993
rect 570 3887 604 3921
rect 642 3887 676 3921
rect 570 3815 604 3849
rect 642 3815 676 3849
rect 570 3743 604 3777
rect 642 3743 676 3777
rect 570 3671 604 3705
rect 642 3671 676 3705
rect 570 3599 604 3633
rect 642 3599 676 3633
rect 570 3527 604 3561
rect 642 3527 676 3561
rect 570 3455 604 3489
rect 642 3455 676 3489
rect 570 3383 604 3417
rect 642 3383 676 3417
rect 570 3311 604 3345
rect 642 3311 676 3345
rect 570 3239 604 3273
rect 642 3239 676 3273
rect 570 3167 604 3201
rect 642 3167 676 3201
rect 570 3095 604 3129
rect 642 3095 676 3129
rect 570 3023 604 3057
rect 642 3023 676 3057
rect 570 2951 604 2985
rect 642 2951 676 2985
rect 570 2879 604 2913
rect 642 2879 676 2913
rect 570 2807 604 2841
rect 642 2807 676 2841
rect 570 2735 604 2769
rect 642 2735 676 2769
rect 570 2663 604 2697
rect 642 2663 676 2697
rect 570 2591 604 2625
rect 642 2591 676 2625
rect 570 2519 604 2553
rect 642 2519 676 2553
rect 570 2447 604 2481
rect 642 2447 676 2481
rect 570 2375 604 2409
rect 642 2375 676 2409
rect 570 2303 604 2337
rect 642 2303 676 2337
rect 570 2231 604 2265
rect 642 2231 676 2265
rect 570 2159 604 2193
rect 642 2159 676 2193
rect 570 2087 604 2121
rect 642 2087 676 2121
rect 570 2015 604 2049
rect 642 2015 676 2049
rect 570 1943 604 1977
rect 642 1943 676 1977
rect 570 1871 604 1905
rect 642 1871 676 1905
rect 570 1799 604 1833
rect 642 1799 676 1833
rect 570 1727 604 1761
rect 642 1727 676 1761
rect 570 1655 604 1689
rect 642 1655 676 1689
rect 570 1583 604 1617
rect 642 1583 676 1617
rect 570 1511 604 1545
rect 642 1511 676 1545
rect 570 1439 604 1473
rect 642 1439 676 1473
rect 570 1367 604 1401
rect 642 1367 676 1401
rect 570 1295 604 1329
rect 642 1295 676 1329
rect 570 1223 604 1257
rect 642 1223 676 1257
rect 570 1151 604 1185
rect 642 1151 676 1185
rect 570 1079 604 1113
rect 642 1079 676 1113
rect 570 1007 604 1041
rect 642 1007 676 1041
rect 570 935 604 969
rect 642 935 676 969
rect 570 863 604 897
rect 642 863 676 897
rect 570 791 604 825
rect 642 791 676 825
rect 570 719 604 753
rect 642 719 676 753
rect 570 647 604 681
rect 642 647 676 681
rect 570 575 604 609
rect 642 575 676 609
rect 570 503 604 537
rect 642 503 676 537
rect 570 431 604 465
rect 642 431 676 465
rect 570 359 604 393
rect 642 359 676 393
rect 570 287 604 321
rect 642 287 676 321
rect 570 215 604 249
rect 642 215 676 249
rect 570 143 604 177
rect 642 143 676 177
rect 570 71 604 105
rect 642 71 676 105
<< poly >>
rect 157 6130 557 6146
rect 157 6096 196 6130
rect 230 6096 268 6130
rect 302 6096 340 6130
rect 374 6096 412 6130
rect 446 6096 484 6130
rect 518 6096 557 6130
rect 157 6040 557 6096
rect 157 0 557 40
<< polycont >>
rect 196 6096 230 6130
rect 268 6096 302 6130
rect 340 6096 374 6130
rect 412 6096 446 6130
rect 484 6096 518 6130
<< locali >>
rect 180 6096 196 6130
rect 230 6096 268 6130
rect 302 6096 340 6130
rect 374 6096 412 6130
rect 446 6096 484 6130
rect 518 6096 534 6130
rect 38 6009 144 6025
rect 38 55 144 71
rect 570 6009 676 6025
rect 570 55 676 71
<< viali >>
rect 196 6096 230 6130
rect 268 6096 302 6130
rect 340 6096 374 6130
rect 412 6096 446 6130
rect 484 6096 518 6130
rect 38 5975 72 6009
rect 72 5975 110 6009
rect 110 5975 144 6009
rect 38 5937 144 5975
rect 38 5903 72 5937
rect 72 5903 110 5937
rect 110 5903 144 5937
rect 38 5865 144 5903
rect 38 5831 72 5865
rect 72 5831 110 5865
rect 110 5831 144 5865
rect 38 5793 144 5831
rect 38 5759 72 5793
rect 72 5759 110 5793
rect 110 5759 144 5793
rect 38 5721 144 5759
rect 38 5687 72 5721
rect 72 5687 110 5721
rect 110 5687 144 5721
rect 38 5649 144 5687
rect 38 5615 72 5649
rect 72 5615 110 5649
rect 110 5615 144 5649
rect 38 5577 144 5615
rect 38 5543 72 5577
rect 72 5543 110 5577
rect 110 5543 144 5577
rect 38 5505 144 5543
rect 38 5471 72 5505
rect 72 5471 110 5505
rect 110 5471 144 5505
rect 38 5433 144 5471
rect 38 5399 72 5433
rect 72 5399 110 5433
rect 110 5399 144 5433
rect 38 5361 144 5399
rect 38 5327 72 5361
rect 72 5327 110 5361
rect 110 5327 144 5361
rect 38 5289 144 5327
rect 38 5255 72 5289
rect 72 5255 110 5289
rect 110 5255 144 5289
rect 38 5217 144 5255
rect 38 5183 72 5217
rect 72 5183 110 5217
rect 110 5183 144 5217
rect 38 5145 144 5183
rect 38 5111 72 5145
rect 72 5111 110 5145
rect 110 5111 144 5145
rect 38 5073 144 5111
rect 38 5039 72 5073
rect 72 5039 110 5073
rect 110 5039 144 5073
rect 38 5001 144 5039
rect 38 4967 72 5001
rect 72 4967 110 5001
rect 110 4967 144 5001
rect 38 4929 144 4967
rect 38 4895 72 4929
rect 72 4895 110 4929
rect 110 4895 144 4929
rect 38 4857 144 4895
rect 38 4823 72 4857
rect 72 4823 110 4857
rect 110 4823 144 4857
rect 38 4785 144 4823
rect 38 4751 72 4785
rect 72 4751 110 4785
rect 110 4751 144 4785
rect 38 4713 144 4751
rect 38 4679 72 4713
rect 72 4679 110 4713
rect 110 4679 144 4713
rect 38 4641 144 4679
rect 38 4607 72 4641
rect 72 4607 110 4641
rect 110 4607 144 4641
rect 38 4569 144 4607
rect 38 4535 72 4569
rect 72 4535 110 4569
rect 110 4535 144 4569
rect 38 4497 144 4535
rect 38 4463 72 4497
rect 72 4463 110 4497
rect 110 4463 144 4497
rect 38 4425 144 4463
rect 38 4391 72 4425
rect 72 4391 110 4425
rect 110 4391 144 4425
rect 38 4353 144 4391
rect 38 4319 72 4353
rect 72 4319 110 4353
rect 110 4319 144 4353
rect 38 4281 144 4319
rect 38 4247 72 4281
rect 72 4247 110 4281
rect 110 4247 144 4281
rect 38 4209 144 4247
rect 38 4175 72 4209
rect 72 4175 110 4209
rect 110 4175 144 4209
rect 38 4137 144 4175
rect 38 4103 72 4137
rect 72 4103 110 4137
rect 110 4103 144 4137
rect 38 4065 144 4103
rect 38 4031 72 4065
rect 72 4031 110 4065
rect 110 4031 144 4065
rect 38 3993 144 4031
rect 38 3959 72 3993
rect 72 3959 110 3993
rect 110 3959 144 3993
rect 38 3921 144 3959
rect 38 3887 72 3921
rect 72 3887 110 3921
rect 110 3887 144 3921
rect 38 3849 144 3887
rect 38 3815 72 3849
rect 72 3815 110 3849
rect 110 3815 144 3849
rect 38 3777 144 3815
rect 38 3743 72 3777
rect 72 3743 110 3777
rect 110 3743 144 3777
rect 38 3705 144 3743
rect 38 3671 72 3705
rect 72 3671 110 3705
rect 110 3671 144 3705
rect 38 3633 144 3671
rect 38 3599 72 3633
rect 72 3599 110 3633
rect 110 3599 144 3633
rect 38 3561 144 3599
rect 38 3527 72 3561
rect 72 3527 110 3561
rect 110 3527 144 3561
rect 38 3489 144 3527
rect 38 3455 72 3489
rect 72 3455 110 3489
rect 110 3455 144 3489
rect 38 3417 144 3455
rect 38 3383 72 3417
rect 72 3383 110 3417
rect 110 3383 144 3417
rect 38 3345 144 3383
rect 38 3311 72 3345
rect 72 3311 110 3345
rect 110 3311 144 3345
rect 38 3273 144 3311
rect 38 3239 72 3273
rect 72 3239 110 3273
rect 110 3239 144 3273
rect 38 3201 144 3239
rect 38 3167 72 3201
rect 72 3167 110 3201
rect 110 3167 144 3201
rect 38 3129 144 3167
rect 38 3095 72 3129
rect 72 3095 110 3129
rect 110 3095 144 3129
rect 38 3057 144 3095
rect 38 3023 72 3057
rect 72 3023 110 3057
rect 110 3023 144 3057
rect 38 2985 144 3023
rect 38 2951 72 2985
rect 72 2951 110 2985
rect 110 2951 144 2985
rect 38 2913 144 2951
rect 38 2879 72 2913
rect 72 2879 110 2913
rect 110 2879 144 2913
rect 38 2841 144 2879
rect 38 2807 72 2841
rect 72 2807 110 2841
rect 110 2807 144 2841
rect 38 2769 144 2807
rect 38 2735 72 2769
rect 72 2735 110 2769
rect 110 2735 144 2769
rect 38 2697 144 2735
rect 38 2663 72 2697
rect 72 2663 110 2697
rect 110 2663 144 2697
rect 38 2625 144 2663
rect 38 2591 72 2625
rect 72 2591 110 2625
rect 110 2591 144 2625
rect 38 2553 144 2591
rect 38 2519 72 2553
rect 72 2519 110 2553
rect 110 2519 144 2553
rect 38 2481 144 2519
rect 38 2447 72 2481
rect 72 2447 110 2481
rect 110 2447 144 2481
rect 38 2409 144 2447
rect 38 2375 72 2409
rect 72 2375 110 2409
rect 110 2375 144 2409
rect 38 2337 144 2375
rect 38 2303 72 2337
rect 72 2303 110 2337
rect 110 2303 144 2337
rect 38 2265 144 2303
rect 38 2231 72 2265
rect 72 2231 110 2265
rect 110 2231 144 2265
rect 38 2193 144 2231
rect 38 2159 72 2193
rect 72 2159 110 2193
rect 110 2159 144 2193
rect 38 2121 144 2159
rect 38 2087 72 2121
rect 72 2087 110 2121
rect 110 2087 144 2121
rect 38 2049 144 2087
rect 38 2015 72 2049
rect 72 2015 110 2049
rect 110 2015 144 2049
rect 38 1977 144 2015
rect 38 1943 72 1977
rect 72 1943 110 1977
rect 110 1943 144 1977
rect 38 1905 144 1943
rect 38 1871 72 1905
rect 72 1871 110 1905
rect 110 1871 144 1905
rect 38 1833 144 1871
rect 38 1799 72 1833
rect 72 1799 110 1833
rect 110 1799 144 1833
rect 38 1761 144 1799
rect 38 1727 72 1761
rect 72 1727 110 1761
rect 110 1727 144 1761
rect 38 1689 144 1727
rect 38 1655 72 1689
rect 72 1655 110 1689
rect 110 1655 144 1689
rect 38 1617 144 1655
rect 38 1583 72 1617
rect 72 1583 110 1617
rect 110 1583 144 1617
rect 38 1545 144 1583
rect 38 1511 72 1545
rect 72 1511 110 1545
rect 110 1511 144 1545
rect 38 1473 144 1511
rect 38 1439 72 1473
rect 72 1439 110 1473
rect 110 1439 144 1473
rect 38 1401 144 1439
rect 38 1367 72 1401
rect 72 1367 110 1401
rect 110 1367 144 1401
rect 38 1329 144 1367
rect 38 1295 72 1329
rect 72 1295 110 1329
rect 110 1295 144 1329
rect 38 1257 144 1295
rect 38 1223 72 1257
rect 72 1223 110 1257
rect 110 1223 144 1257
rect 38 1185 144 1223
rect 38 1151 72 1185
rect 72 1151 110 1185
rect 110 1151 144 1185
rect 38 1113 144 1151
rect 38 1079 72 1113
rect 72 1079 110 1113
rect 110 1079 144 1113
rect 38 1041 144 1079
rect 38 1007 72 1041
rect 72 1007 110 1041
rect 110 1007 144 1041
rect 38 969 144 1007
rect 38 935 72 969
rect 72 935 110 969
rect 110 935 144 969
rect 38 897 144 935
rect 38 863 72 897
rect 72 863 110 897
rect 110 863 144 897
rect 38 825 144 863
rect 38 791 72 825
rect 72 791 110 825
rect 110 791 144 825
rect 38 753 144 791
rect 38 719 72 753
rect 72 719 110 753
rect 110 719 144 753
rect 38 681 144 719
rect 38 647 72 681
rect 72 647 110 681
rect 110 647 144 681
rect 38 609 144 647
rect 38 575 72 609
rect 72 575 110 609
rect 110 575 144 609
rect 38 537 144 575
rect 38 503 72 537
rect 72 503 110 537
rect 110 503 144 537
rect 38 465 144 503
rect 38 431 72 465
rect 72 431 110 465
rect 110 431 144 465
rect 38 393 144 431
rect 38 359 72 393
rect 72 359 110 393
rect 110 359 144 393
rect 38 321 144 359
rect 38 287 72 321
rect 72 287 110 321
rect 110 287 144 321
rect 38 249 144 287
rect 38 215 72 249
rect 72 215 110 249
rect 110 215 144 249
rect 38 177 144 215
rect 38 143 72 177
rect 72 143 110 177
rect 110 143 144 177
rect 38 105 144 143
rect 38 71 72 105
rect 72 71 110 105
rect 110 71 144 105
rect 570 5975 604 6009
rect 604 5975 642 6009
rect 642 5975 676 6009
rect 570 5937 676 5975
rect 570 5903 604 5937
rect 604 5903 642 5937
rect 642 5903 676 5937
rect 570 5865 676 5903
rect 570 5831 604 5865
rect 604 5831 642 5865
rect 642 5831 676 5865
rect 570 5793 676 5831
rect 570 5759 604 5793
rect 604 5759 642 5793
rect 642 5759 676 5793
rect 570 5721 676 5759
rect 570 5687 604 5721
rect 604 5687 642 5721
rect 642 5687 676 5721
rect 570 5649 676 5687
rect 570 5615 604 5649
rect 604 5615 642 5649
rect 642 5615 676 5649
rect 570 5577 676 5615
rect 570 5543 604 5577
rect 604 5543 642 5577
rect 642 5543 676 5577
rect 570 5505 676 5543
rect 570 5471 604 5505
rect 604 5471 642 5505
rect 642 5471 676 5505
rect 570 5433 676 5471
rect 570 5399 604 5433
rect 604 5399 642 5433
rect 642 5399 676 5433
rect 570 5361 676 5399
rect 570 5327 604 5361
rect 604 5327 642 5361
rect 642 5327 676 5361
rect 570 5289 676 5327
rect 570 5255 604 5289
rect 604 5255 642 5289
rect 642 5255 676 5289
rect 570 5217 676 5255
rect 570 5183 604 5217
rect 604 5183 642 5217
rect 642 5183 676 5217
rect 570 5145 676 5183
rect 570 5111 604 5145
rect 604 5111 642 5145
rect 642 5111 676 5145
rect 570 5073 676 5111
rect 570 5039 604 5073
rect 604 5039 642 5073
rect 642 5039 676 5073
rect 570 5001 676 5039
rect 570 4967 604 5001
rect 604 4967 642 5001
rect 642 4967 676 5001
rect 570 4929 676 4967
rect 570 4895 604 4929
rect 604 4895 642 4929
rect 642 4895 676 4929
rect 570 4857 676 4895
rect 570 4823 604 4857
rect 604 4823 642 4857
rect 642 4823 676 4857
rect 570 4785 676 4823
rect 570 4751 604 4785
rect 604 4751 642 4785
rect 642 4751 676 4785
rect 570 4713 676 4751
rect 570 4679 604 4713
rect 604 4679 642 4713
rect 642 4679 676 4713
rect 570 4641 676 4679
rect 570 4607 604 4641
rect 604 4607 642 4641
rect 642 4607 676 4641
rect 570 4569 676 4607
rect 570 4535 604 4569
rect 604 4535 642 4569
rect 642 4535 676 4569
rect 570 4497 676 4535
rect 570 4463 604 4497
rect 604 4463 642 4497
rect 642 4463 676 4497
rect 570 4425 676 4463
rect 570 4391 604 4425
rect 604 4391 642 4425
rect 642 4391 676 4425
rect 570 4353 676 4391
rect 570 4319 604 4353
rect 604 4319 642 4353
rect 642 4319 676 4353
rect 570 4281 676 4319
rect 570 4247 604 4281
rect 604 4247 642 4281
rect 642 4247 676 4281
rect 570 4209 676 4247
rect 570 4175 604 4209
rect 604 4175 642 4209
rect 642 4175 676 4209
rect 570 4137 676 4175
rect 570 4103 604 4137
rect 604 4103 642 4137
rect 642 4103 676 4137
rect 570 4065 676 4103
rect 570 4031 604 4065
rect 604 4031 642 4065
rect 642 4031 676 4065
rect 570 3993 676 4031
rect 570 3959 604 3993
rect 604 3959 642 3993
rect 642 3959 676 3993
rect 570 3921 676 3959
rect 570 3887 604 3921
rect 604 3887 642 3921
rect 642 3887 676 3921
rect 570 3849 676 3887
rect 570 3815 604 3849
rect 604 3815 642 3849
rect 642 3815 676 3849
rect 570 3777 676 3815
rect 570 3743 604 3777
rect 604 3743 642 3777
rect 642 3743 676 3777
rect 570 3705 676 3743
rect 570 3671 604 3705
rect 604 3671 642 3705
rect 642 3671 676 3705
rect 570 3633 676 3671
rect 570 3599 604 3633
rect 604 3599 642 3633
rect 642 3599 676 3633
rect 570 3561 676 3599
rect 570 3527 604 3561
rect 604 3527 642 3561
rect 642 3527 676 3561
rect 570 3489 676 3527
rect 570 3455 604 3489
rect 604 3455 642 3489
rect 642 3455 676 3489
rect 570 3417 676 3455
rect 570 3383 604 3417
rect 604 3383 642 3417
rect 642 3383 676 3417
rect 570 3345 676 3383
rect 570 3311 604 3345
rect 604 3311 642 3345
rect 642 3311 676 3345
rect 570 3273 676 3311
rect 570 3239 604 3273
rect 604 3239 642 3273
rect 642 3239 676 3273
rect 570 3201 676 3239
rect 570 3167 604 3201
rect 604 3167 642 3201
rect 642 3167 676 3201
rect 570 3129 676 3167
rect 570 3095 604 3129
rect 604 3095 642 3129
rect 642 3095 676 3129
rect 570 3057 676 3095
rect 570 3023 604 3057
rect 604 3023 642 3057
rect 642 3023 676 3057
rect 570 2985 676 3023
rect 570 2951 604 2985
rect 604 2951 642 2985
rect 642 2951 676 2985
rect 570 2913 676 2951
rect 570 2879 604 2913
rect 604 2879 642 2913
rect 642 2879 676 2913
rect 570 2841 676 2879
rect 570 2807 604 2841
rect 604 2807 642 2841
rect 642 2807 676 2841
rect 570 2769 676 2807
rect 570 2735 604 2769
rect 604 2735 642 2769
rect 642 2735 676 2769
rect 570 2697 676 2735
rect 570 2663 604 2697
rect 604 2663 642 2697
rect 642 2663 676 2697
rect 570 2625 676 2663
rect 570 2591 604 2625
rect 604 2591 642 2625
rect 642 2591 676 2625
rect 570 2553 676 2591
rect 570 2519 604 2553
rect 604 2519 642 2553
rect 642 2519 676 2553
rect 570 2481 676 2519
rect 570 2447 604 2481
rect 604 2447 642 2481
rect 642 2447 676 2481
rect 570 2409 676 2447
rect 570 2375 604 2409
rect 604 2375 642 2409
rect 642 2375 676 2409
rect 570 2337 676 2375
rect 570 2303 604 2337
rect 604 2303 642 2337
rect 642 2303 676 2337
rect 570 2265 676 2303
rect 570 2231 604 2265
rect 604 2231 642 2265
rect 642 2231 676 2265
rect 570 2193 676 2231
rect 570 2159 604 2193
rect 604 2159 642 2193
rect 642 2159 676 2193
rect 570 2121 676 2159
rect 570 2087 604 2121
rect 604 2087 642 2121
rect 642 2087 676 2121
rect 570 2049 676 2087
rect 570 2015 604 2049
rect 604 2015 642 2049
rect 642 2015 676 2049
rect 570 1977 676 2015
rect 570 1943 604 1977
rect 604 1943 642 1977
rect 642 1943 676 1977
rect 570 1905 676 1943
rect 570 1871 604 1905
rect 604 1871 642 1905
rect 642 1871 676 1905
rect 570 1833 676 1871
rect 570 1799 604 1833
rect 604 1799 642 1833
rect 642 1799 676 1833
rect 570 1761 676 1799
rect 570 1727 604 1761
rect 604 1727 642 1761
rect 642 1727 676 1761
rect 570 1689 676 1727
rect 570 1655 604 1689
rect 604 1655 642 1689
rect 642 1655 676 1689
rect 570 1617 676 1655
rect 570 1583 604 1617
rect 604 1583 642 1617
rect 642 1583 676 1617
rect 570 1545 676 1583
rect 570 1511 604 1545
rect 604 1511 642 1545
rect 642 1511 676 1545
rect 570 1473 676 1511
rect 570 1439 604 1473
rect 604 1439 642 1473
rect 642 1439 676 1473
rect 570 1401 676 1439
rect 570 1367 604 1401
rect 604 1367 642 1401
rect 642 1367 676 1401
rect 570 1329 676 1367
rect 570 1295 604 1329
rect 604 1295 642 1329
rect 642 1295 676 1329
rect 570 1257 676 1295
rect 570 1223 604 1257
rect 604 1223 642 1257
rect 642 1223 676 1257
rect 570 1185 676 1223
rect 570 1151 604 1185
rect 604 1151 642 1185
rect 642 1151 676 1185
rect 570 1113 676 1151
rect 570 1079 604 1113
rect 604 1079 642 1113
rect 642 1079 676 1113
rect 570 1041 676 1079
rect 570 1007 604 1041
rect 604 1007 642 1041
rect 642 1007 676 1041
rect 570 969 676 1007
rect 570 935 604 969
rect 604 935 642 969
rect 642 935 676 969
rect 570 897 676 935
rect 570 863 604 897
rect 604 863 642 897
rect 642 863 676 897
rect 570 825 676 863
rect 570 791 604 825
rect 604 791 642 825
rect 642 791 676 825
rect 570 753 676 791
rect 570 719 604 753
rect 604 719 642 753
rect 642 719 676 753
rect 570 681 676 719
rect 570 647 604 681
rect 604 647 642 681
rect 642 647 676 681
rect 570 609 676 647
rect 570 575 604 609
rect 604 575 642 609
rect 642 575 676 609
rect 570 537 676 575
rect 570 503 604 537
rect 604 503 642 537
rect 642 503 676 537
rect 570 465 676 503
rect 570 431 604 465
rect 604 431 642 465
rect 642 431 676 465
rect 570 393 676 431
rect 570 359 604 393
rect 604 359 642 393
rect 642 359 676 393
rect 570 321 676 359
rect 570 287 604 321
rect 604 287 642 321
rect 642 287 676 321
rect 570 249 676 287
rect 570 215 604 249
rect 604 215 642 249
rect 642 215 676 249
rect 570 177 676 215
rect 570 143 604 177
rect 604 143 642 177
rect 642 143 676 177
rect 570 105 676 143
rect 570 71 604 105
rect 604 71 642 105
rect 642 71 676 105
<< metal1 >>
rect 184 6130 530 6136
rect 184 6096 196 6130
rect 230 6096 268 6130
rect 302 6096 340 6130
rect 374 6096 412 6130
rect 446 6096 484 6130
rect 518 6096 530 6130
rect 184 6090 530 6096
rect 32 6009 150 6021
rect 32 71 38 6009
rect 144 71 150 6009
rect 32 59 150 71
rect 564 6009 682 6021
rect 564 71 570 6009
rect 676 71 682 6009
rect 564 59 682 71
<< end >>
