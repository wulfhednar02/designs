magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -5 0 375 2592
<< l68d20 >>
rect 0 0 370 720
<< l68d44 >>
rect 110 460 260 610
rect 110 110 260 260
<< l69d20 >>
rect -5 0 375 1495
<< l70d44 >>
rect 85 1610 285 1810
rect 85 2010 285 2210
<< l69d44 >>
rect 85 1210 285 1410
rect 85 810 285 1010
<< l71d20 >>
rect -5 1520 375 2300
rect 35 2300 335 2592
<< l70d20 >>
rect -5 720 375 2300
<< end >>
