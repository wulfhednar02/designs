magic
tech sky130A
timestamp 1699066547
<< end >>
