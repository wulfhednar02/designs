magic
tech sky130A
magscale 1 2
timestamp 1698982078
<< metal1 >>
rect 1 133 75 144
rect 1 81 12 133
rect 64 81 75 133
rect 1 63 75 81
rect 1 11 12 63
rect 64 11 75 63
rect 1 0 75 11
<< via1 >>
rect 12 81 64 133
rect 12 11 64 63
<< metal2 >>
rect 0 290 76 298
rect 0 234 10 290
rect 66 234 76 290
rect 0 210 76 234
rect 0 154 10 210
rect 66 154 76 210
rect 0 133 76 154
rect 0 81 12 133
rect 64 81 76 133
rect 0 63 76 81
rect 0 11 12 63
rect 64 11 76 63
rect 0 0 76 11
<< via2 >>
rect 10 234 66 290
rect 10 154 66 210
<< metal3 >>
rect 0 294 76 299
rect 0 230 6 294
rect 70 230 76 294
rect 0 214 76 230
rect 0 150 6 214
rect 70 150 76 214
rect 0 144 76 150
<< via3 >>
rect 6 290 70 294
rect 6 234 10 290
rect 10 234 66 290
rect 66 234 70 290
rect 6 230 70 234
rect 6 210 70 214
rect 6 154 10 210
rect 10 154 66 210
rect 66 154 70 210
rect 6 150 70 154
<< metal4 >>
rect 8 299 68 518
rect 0 294 76 299
rect 0 230 6 294
rect 70 230 76 294
rect 0 214 76 230
rect 0 150 6 214
rect 70 150 76 214
rect 0 144 76 150
<< end >>
