magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -190 -240 10310 2960
<< l66d20 >>
rect 395 105 545 1025
rect 815 105 965 1025
rect 1235 105 1385 1025
rect 1655 105 1805 1025
rect 2075 105 2225 1025
rect 2495 105 2645 1025
rect 395 1025 2645 1295
rect 395 1295 545 2615
rect 815 1295 965 2615
rect 1235 1295 1385 2615
rect 1655 1295 1805 2615
rect 2075 1295 2225 2615
rect 2495 1295 2645 2615
rect 2915 105 3065 1025
rect 3335 105 3485 1025
rect 3755 105 3905 1025
rect 4175 105 4325 1025
rect 4595 105 4745 1025
rect 5015 105 5165 1025
rect 5435 105 5585 1025
rect 5855 105 6005 1025
rect 6275 105 6425 1025
rect 6695 105 6845 1025
rect 7115 105 7265 1025
rect 7535 105 7685 1025
rect 7955 105 8105 1025
rect 8375 105 8525 1025
rect 8795 105 8945 1025
rect 9215 105 9365 1025
rect 2915 1025 9385 1295
rect 2915 1295 3065 2615
rect 3335 1295 3485 2615
rect 3755 1295 3905 2615
rect 4175 1295 4325 2615
rect 4595 1295 4745 2615
rect 5015 1295 5165 2615
rect 5435 1295 5585 2615
rect 5855 1295 6005 2615
rect 6275 1295 6425 2615
rect 6695 1295 6845 2615
rect 7115 1295 7265 2615
rect 7535 1295 7685 2615
rect 7955 1295 8105 2615
rect 8375 1295 8525 2615
rect 8795 1295 8945 2615
rect 9215 1295 9365 2615
<< l94d20 >>
rect 0 1355 10120 2910
<< l66d44 >>
rect 4715 1075 4885 1245
rect 4795 2225 4965 2395
rect 4795 1885 4965 2055
rect 4795 1545 4965 1715
rect 4795 655 4965 825
rect 4795 315 4965 485
rect 5055 1075 5225 1245
rect 5215 2255 5385 2425
rect 5215 1915 5385 2085
rect 5215 315 5385 485
rect 5395 1075 5565 1245
rect 5635 2225 5805 2395
rect 5635 1885 5805 2055
rect 5635 1545 5805 1715
rect 5635 655 5805 825
rect 5635 315 5805 485
rect 5735 1075 5905 1245
rect 6055 2255 6225 2425
rect 6055 1915 6225 2085
rect 6055 315 6225 485
rect 6075 1075 6245 1245
rect 6415 1075 6585 1245
rect 6475 2225 6645 2395
rect 6475 1885 6645 2055
rect 6475 1545 6645 1715
rect 6475 655 6645 825
rect 6475 315 6645 485
rect 6755 1075 6925 1245
rect 6895 2255 7065 2425
rect 6895 1915 7065 2085
rect 9415 315 9585 485
rect 6895 315 7065 485
rect 7095 1075 7265 1245
rect 7315 2225 7485 2395
rect 7315 1885 7485 2055
rect 7315 1545 7485 1715
rect 7315 655 7485 825
rect 7315 315 7485 485
rect 7435 1075 7605 1245
rect 7735 2255 7905 2425
rect 7735 1915 7905 2085
rect 7735 315 7905 485
rect 7775 1075 7945 1245
rect 8115 1075 8285 1245
rect 8155 2225 8325 2395
rect 8155 1885 8325 2055
rect 8155 1545 8325 1715
rect 8155 655 8325 825
rect 8155 315 8325 485
rect 8455 1075 8625 1245
rect 8575 2255 8745 2425
rect 8575 1915 8745 2085
rect 8575 315 8745 485
rect 8795 1075 8965 1245
rect 8995 2225 9165 2395
rect 8995 1885 9165 2055
rect 8995 1545 9165 1715
rect 8995 655 9165 825
rect 8995 315 9165 485
rect 9135 1075 9305 1245
rect 9415 2255 9585 2425
rect 9415 1915 9585 2085
rect 1015 1915 1185 2085
rect 1015 315 1185 485
rect 1195 1075 1365 1245
rect 1435 2225 1605 2395
rect 1855 1915 2025 2085
rect 1855 315 2025 485
rect 1875 1075 2045 1245
rect 2215 1075 2385 1245
rect 2275 2225 2445 2395
rect 2275 1885 2445 2055
rect 2275 1545 2445 1715
rect 2275 655 2445 825
rect 2275 315 2445 485
rect 2695 2255 2865 2425
rect 3955 1885 4125 2055
rect 3955 1545 4125 1715
rect 3955 655 4125 825
rect 3955 315 4125 485
rect 4035 1075 4205 1245
rect 4375 2255 4545 2425
rect 4375 1915 4545 2085
rect 4375 1075 4545 1245
rect 4375 315 4545 485
rect 1435 1885 1605 2055
rect 1435 1545 1605 1715
rect 1435 655 1605 825
rect 1435 315 1605 485
rect 1535 1075 1705 1245
rect 1855 2255 2025 2425
rect 595 1885 765 2055
rect 595 1545 765 1715
rect 595 655 765 825
rect 595 315 765 485
rect 855 1075 1025 1245
rect 1015 2255 1185 2425
rect 175 2255 345 2425
rect 175 1915 345 2085
rect 175 1575 345 1745
rect 175 655 345 825
rect 175 315 345 485
rect 515 1075 685 1245
rect 595 2225 765 2395
rect 3535 2255 3705 2425
rect 3535 1915 3705 2085
rect 3535 315 3705 485
rect 3695 1075 3865 1245
rect 3955 2225 4125 2395
rect 2695 1915 2865 2085
rect 2695 315 2865 485
rect 3015 1075 3185 1245
rect 3115 2225 3285 2395
rect 3115 1885 3285 2055
rect 3115 1545 3285 1715
rect 3115 655 3285 825
rect 3115 315 3285 485
rect 3355 1075 3525 1245
<< l67d44 >>
rect 8425 2635 8595 2805
rect 8425 -85 8595 85
rect 145 2635 315 2805
rect 145 -85 315 85
rect 605 2635 775 2805
rect 605 -85 775 85
rect 1065 2635 1235 2805
rect 1065 -85 1235 85
rect 1525 2635 1695 2805
rect 1525 -85 1695 85
rect 1985 2635 2155 2805
rect 1985 -85 2155 85
rect 2445 2635 2615 2805
rect 2445 -85 2615 85
rect 2905 2635 3075 2805
rect 2905 -85 3075 85
rect 3365 2635 3535 2805
rect 3365 -85 3535 85
rect 3825 2635 3995 2805
rect 3825 -85 3995 85
rect 4285 2635 4455 2805
rect 4285 -85 4455 85
rect 4745 2635 4915 2805
rect 4745 -85 4915 85
rect 5205 2635 5375 2805
rect 5205 -85 5375 85
rect 5665 2635 5835 2805
rect 5665 -85 5835 85
rect 6125 2635 6295 2805
rect 6125 -85 6295 85
rect 6585 2635 6755 2805
rect 6585 -85 6755 85
rect 7045 2635 7215 2805
rect 7045 -85 7215 85
rect 7505 2635 7675 2805
rect 7505 -85 7675 85
rect 7965 2635 8135 2805
rect 7965 -85 8135 85
rect 8885 2635 9055 2805
rect 8885 -85 9055 85
rect 9345 2635 9515 2805
rect 9345 -85 9515 85
rect 9805 2635 9975 2805
rect 9805 -85 9975 85
<< l95d20 >>
rect 0 975 10120 1345
<< l67d20 >>
rect 0 -85 10120 85
rect 1015 85 1185 565
rect 1855 85 2025 565
rect 2695 85 2865 565
rect 3535 85 3705 565
rect 4375 85 4545 565
rect 5215 85 5385 565
rect 6055 85 6225 565
rect 6895 85 7065 565
rect 7735 85 7905 565
rect 8575 85 8745 565
rect 9415 85 9585 565
rect 175 85 345 905
rect 175 1445 345 2635
rect 1015 1835 1185 2635
rect 1855 1835 2025 2635
rect 2695 1835 2865 2635
rect 3535 1835 3705 2635
rect 4375 1835 4545 2635
rect 5215 1835 5385 2635
rect 6055 1835 6225 2635
rect 6895 1835 7065 2635
rect 7735 1835 7905 2635
rect 8575 1835 8745 2635
rect 9415 1835 9585 2635
rect 0 2635 10120 2805
rect 515 260 845 735
rect 1355 260 1685 735
rect 2195 260 2525 735
rect 515 735 2865 905
rect 2690 905 2865 1075
rect 2690 1075 9410 1275
rect 2690 1275 2865 1445
rect 515 1445 2865 1615
rect 515 1615 845 2465
rect 1355 1615 1685 2465
rect 2195 1615 2525 2465
rect 3035 255 3285 260
rect 3955 255 4125 260
rect 4795 255 4965 260
rect 3035 260 3365 735
rect 3875 260 4205 735
rect 4715 260 5045 735
rect 5555 260 5885 735
rect 6395 260 6725 735
rect 7235 260 7565 735
rect 8075 260 8405 735
rect 8915 260 9245 735
rect 9760 365 10035 735
rect 3035 735 10035 905
rect 9655 905 10035 1445
rect 3035 1445 10035 1615
rect 9760 1615 10035 2360
rect 3035 1615 3365 2465
rect 3875 1615 4205 2465
rect 4715 1615 5045 2465
rect 5555 1615 5885 2465
rect 6395 1615 6725 2465
rect 7235 1615 7565 2465
rect 8075 1615 8405 2465
rect 8915 1615 9245 2465
rect 85 1075 2485 1275
<< l68d20 >>
rect 0 -240 10120 240
rect 0 2480 10120 2960
<< l65d20 >>
rect 135 1485 9625 2485
rect 135 235 9625 885
<< l93d44 >>
rect 0 -190 10120 1015
<< l64d20 >>
rect -190 1305 10310 2910
<< l68d16 >>
rect 150 -85 320 85
rect 150 2635 320 2805
<< l236d0 >>
rect 0 0 10120 2720
<< l122d16 >>
rect 150 -85 320 85
<< l64d16 >>
rect 150 2635 320 2805
<< l81d4 >>
rect 0 0 10120 2720
<< l78d44 >>
rect 0 1250 10120 2720
<< l67d16 >>
rect 1530 1105 1700 1275
rect 1990 1105 2160 1275
rect 9805 1445 9975 1615
rect 9805 1105 9975 1275
<< labels >>
rlabel l67d5 2075 1190 2075 1190 0 A
rlabel l67d5 1615 1190 1615 1190 0 A
rlabel l67d5 9890 1190 9890 1190 0 X
rlabel l67d5 9890 1530 9890 1530 0 X
rlabel l64d59 235 0 235 0 0 VNB
rlabel l64d5 235 2720 235 2720 0 VPB
rlabel l68d5 230 0 230 0 0 VGND
rlabel l68d5 230 2720 230 2720 0 VPWR
rlabel l83d44 0 0 0 0 0 buf_16
<< end >>
