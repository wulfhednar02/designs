magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< error_p >>
rect -105 22 -36 91
rect -35 22 35 49
rect 36 22 105 91
rect -105 21 105 22
rect -467 20 34 21
rect 35 20 467 21
rect -467 -21 -36 -20
rect -35 -21 34 -20
rect 36 -21 467 -20
<< xpolycontact >>
rect -36 21 36 458
rect -36 20 -35 21
rect -36 -21 -35 -20
rect 35 20 36 21
rect 35 -21 36 -20
rect -36 -458 36 -21
<< ppolyres >>
rect -35 -21 35 21
<< locali >>
rect -35 20 35 21
rect -35 -21 35 -20
<< viali >>
rect -17 404 17 438
rect -17 332 17 366
rect -17 260 17 294
rect -17 188 17 222
rect -17 116 17 150
rect -17 44 17 78
rect -17 -77 17 -43
rect -17 -149 17 -115
rect -17 -221 17 -187
rect -17 -293 17 -259
rect -17 -365 17 -331
rect -17 -437 17 -403
<< metal1 >>
rect -25 438 25 451
rect -25 404 -17 438
rect 17 404 25 438
rect -25 366 25 404
rect -25 332 -17 366
rect 17 332 25 366
rect -25 294 25 332
rect -25 260 -17 294
rect 17 260 25 294
rect -25 222 25 260
rect -25 188 -17 222
rect 17 188 25 222
rect -25 150 25 188
rect -25 116 -17 150
rect 17 116 25 150
rect -25 78 25 116
rect -25 44 -17 78
rect 17 44 25 78
rect -25 30 25 44
rect -25 -43 25 -30
rect -25 -77 -17 -43
rect 17 -77 25 -43
rect -25 -115 25 -77
rect -25 -149 -17 -115
rect 17 -149 25 -115
rect -25 -187 25 -149
rect -25 -221 -17 -187
rect 17 -221 25 -187
rect -25 -259 25 -221
rect -25 -293 -17 -259
rect 17 -293 25 -259
rect -25 -331 25 -293
rect -25 -365 -17 -331
rect 17 -365 25 -331
rect -25 -403 25 -365
rect -25 -437 -17 -403
rect 17 -437 25 -403
rect -25 -451 25 -437
<< end >>
