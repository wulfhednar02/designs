magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -635 -2485 635 2485
<< l66d20 >>
rect -175 -2285 175 2285
<< l94d20 >>
rect -285 -2395 285 2395
<< l86d20 >>
rect -635 -2485 635 2485
<< l66d44 >>
rect -95 205 95 2205
rect -95 -2205 95 -205
<< l67d44 >>
rect -85 220 85 390
rect -85 580 85 750
rect -85 940 85 1110
rect -85 1300 85 1470
rect -85 1660 85 1830
rect -85 2020 85 2190
rect -85 -2185 85 -2015
rect -85 -1825 85 -1655
rect -85 -1465 85 -1295
rect -85 -1105 85 -935
rect -85 -745 85 -575
rect -85 -385 85 -215
<< l95d20 >>
rect -270 -2380 270 2380
<< l67d20 >>
rect -175 125 175 2285
rect -175 -2285 175 -125
<< l66d13 >>
rect -175 -185 175 185
<< l68d20 >>
rect -125 151 125 2255
rect -125 -2255 125 -151
<< end >>
