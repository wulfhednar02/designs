magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect -125 -200 3445 30540
<< l66d20 >>
rect 660 -200 2660 30200
rect 660 30200 2660 30530
<< l66d44 >>
rect 65 15275 235 15445
rect 425 15275 595 15445
rect 2725 15275 2895 15445
rect 3085 15275 3255 15445
rect 65 22835 235 23005
rect 425 22835 595 23005
rect 2725 22835 2895 23005
rect 3085 22835 3255 23005
rect 65 24275 235 24445
rect 65 24635 235 24805
rect 65 24995 235 25165
rect 65 25355 235 25525
rect 65 25715 235 25885
rect 65 26075 235 26245
rect 65 26435 235 26605
rect 65 26795 235 26965
rect 65 27155 235 27325
rect 65 27515 235 27685
rect 65 27875 235 28045
rect 65 28235 235 28405
rect 65 28595 235 28765
rect 65 28955 235 29125
rect 65 29315 235 29485
rect 65 29675 235 29845
rect 65 23195 235 23365
rect 425 23195 595 23365
rect 425 23555 595 23725
rect 425 23915 595 24085
rect 425 24275 595 24445
rect 425 24635 595 24805
rect 425 24995 595 25165
rect 425 25355 595 25525
rect 425 25715 595 25885
rect 425 26075 595 26245
rect 425 26435 595 26605
rect 425 26795 595 26965
rect 425 27155 595 27325
rect 425 27515 595 27685
rect 425 27875 595 28045
rect 425 28235 595 28405
rect 425 28595 595 28765
rect 425 28955 595 29125
rect 425 29315 595 29485
rect 425 29675 595 29845
rect 65 23555 235 23725
rect 2725 23195 2895 23365
rect 2725 23555 2895 23725
rect 2725 23915 2895 24085
rect 2725 24275 2895 24445
rect 2725 24635 2895 24805
rect 2725 24995 2895 25165
rect 2725 25355 2895 25525
rect 2725 25715 2895 25885
rect 2725 26075 2895 26245
rect 2725 26435 2895 26605
rect 2725 26795 2895 26965
rect 2725 27155 2895 27325
rect 2725 27515 2895 27685
rect 2725 27875 2895 28045
rect 2725 28235 2895 28405
rect 2725 28595 2895 28765
rect 2725 28955 2895 29125
rect 2725 29315 2895 29485
rect 2725 29675 2895 29845
rect 65 23915 235 24085
rect 3085 23195 3255 23365
rect 3085 23555 3255 23725
rect 3085 23915 3255 24085
rect 3085 24275 3255 24445
rect 3085 24635 3255 24805
rect 3085 24995 3255 25165
rect 3085 25355 3255 25525
rect 3085 25715 3255 25885
rect 3085 26075 3255 26245
rect 3085 26435 3255 26605
rect 3085 26795 3255 26965
rect 3085 27155 3255 27325
rect 3085 27515 3255 27685
rect 3085 27875 3255 28045
rect 3085 28235 3255 28405
rect 3085 28595 3255 28765
rect 3085 28955 3255 29125
rect 3085 29315 3255 29485
rect 3085 29675 3255 29845
rect 855 30280 1025 30450
rect 1215 30280 1385 30450
rect 1575 30280 1745 30450
rect 1935 30280 2105 30450
rect 2295 30280 2465 30450
rect 2725 17795 2895 17965
rect 2725 18155 2895 18325
rect 2725 18515 2895 18685
rect 2725 18875 2895 19045
rect 2725 19235 2895 19405
rect 2725 19595 2895 19765
rect 2725 19955 2895 20125
rect 2725 20315 2895 20485
rect 2725 20675 2895 20845
rect 2725 21035 2895 21205
rect 2725 21395 2895 21565
rect 2725 21755 2895 21925
rect 2725 22115 2895 22285
rect 2725 22475 2895 22645
rect 425 16355 595 16525
rect 425 16715 595 16885
rect 425 17075 595 17245
rect 425 17435 595 17605
rect 425 17795 595 17965
rect 425 18155 595 18325
rect 425 18515 595 18685
rect 425 18875 595 19045
rect 425 19235 595 19405
rect 425 19595 595 19765
rect 425 19955 595 20125
rect 425 20315 595 20485
rect 425 20675 595 20845
rect 425 21035 595 21205
rect 425 21395 595 21565
rect 425 21755 595 21925
rect 425 22115 595 22285
rect 425 22475 595 22645
rect 65 17795 235 17965
rect 65 18155 235 18325
rect 65 16355 235 16525
rect 3085 15635 3255 15805
rect 3085 15995 3255 16165
rect 3085 16355 3255 16525
rect 3085 16715 3255 16885
rect 3085 17075 3255 17245
rect 3085 17435 3255 17605
rect 3085 17795 3255 17965
rect 3085 18155 3255 18325
rect 3085 18515 3255 18685
rect 3085 18875 3255 19045
rect 3085 19235 3255 19405
rect 3085 19595 3255 19765
rect 3085 19955 3255 20125
rect 3085 20315 3255 20485
rect 3085 20675 3255 20845
rect 3085 21035 3255 21205
rect 3085 21395 3255 21565
rect 3085 21755 3255 21925
rect 3085 22115 3255 22285
rect 3085 22475 3255 22645
rect 65 18515 235 18685
rect 65 18875 235 19045
rect 65 19235 235 19405
rect 65 19595 235 19765
rect 65 19955 235 20125
rect 65 20315 235 20485
rect 65 20675 235 20845
rect 65 21035 235 21205
rect 65 21395 235 21565
rect 65 21755 235 21925
rect 65 22115 235 22285
rect 65 22475 235 22645
rect 65 16715 235 16885
rect 65 17075 235 17245
rect 65 17435 235 17605
rect 65 15635 235 15805
rect 425 15635 595 15805
rect 425 15995 595 16165
rect 65 15995 235 16165
rect 2725 15635 2895 15805
rect 2725 15995 2895 16165
rect 2725 16355 2895 16525
rect 2725 16715 2895 16885
rect 2725 17075 2895 17245
rect 2725 17435 2895 17605
rect 2725 7715 2895 7885
rect 425 7715 595 7885
rect 3085 7715 3255 7885
rect 65 7715 235 7885
rect 2725 9155 2895 9325
rect 2725 9515 2895 9685
rect 2725 9875 2895 10045
rect 2725 10235 2895 10405
rect 2725 10595 2895 10765
rect 2725 10955 2895 11125
rect 2725 11315 2895 11485
rect 2725 11675 2895 11845
rect 2725 12035 2895 12205
rect 2725 12395 2895 12565
rect 2725 12755 2895 12925
rect 2725 13115 2895 13285
rect 2725 13475 2895 13645
rect 2725 13835 2895 14005
rect 2725 14195 2895 14365
rect 2725 14555 2895 14725
rect 2725 14915 2895 15085
rect 65 14555 235 14725
rect 2725 8075 2895 8245
rect 425 8075 595 8245
rect 425 8435 595 8605
rect 425 8795 595 8965
rect 425 9155 595 9325
rect 425 9515 595 9685
rect 425 9875 595 10045
rect 425 10235 595 10405
rect 425 10595 595 10765
rect 425 10955 595 11125
rect 425 11315 595 11485
rect 425 11675 595 11845
rect 425 12035 595 12205
rect 425 12395 595 12565
rect 425 12755 595 12925
rect 425 13115 595 13285
rect 425 13475 595 13645
rect 425 13835 595 14005
rect 425 14195 595 14365
rect 2725 8435 2895 8605
rect 3085 8075 3255 8245
rect 3085 8435 3255 8605
rect 3085 8795 3255 8965
rect 3085 9155 3255 9325
rect 3085 9515 3255 9685
rect 3085 9875 3255 10045
rect 3085 10235 3255 10405
rect 3085 10595 3255 10765
rect 3085 10955 3255 11125
rect 3085 11315 3255 11485
rect 3085 11675 3255 11845
rect 3085 12035 3255 12205
rect 3085 12395 3255 12565
rect 3085 12755 3255 12925
rect 3085 13115 3255 13285
rect 3085 13475 3255 13645
rect 3085 13835 3255 14005
rect 3085 14195 3255 14365
rect 3085 14555 3255 14725
rect 3085 14915 3255 15085
rect 425 14555 595 14725
rect 425 14915 595 15085
rect 65 14915 235 15085
rect 2725 8795 2895 8965
rect 65 8075 235 8245
rect 65 8435 235 8605
rect 65 8795 235 8965
rect 65 9155 235 9325
rect 65 9515 235 9685
rect 65 9875 235 10045
rect 65 10235 235 10405
rect 65 10595 235 10765
rect 65 10955 235 11125
rect 65 11315 235 11485
rect 65 11675 235 11845
rect 65 12035 235 12205
rect 65 12395 235 12565
rect 65 12755 235 12925
rect 65 13115 235 13285
rect 65 13475 235 13645
rect 65 13835 235 14005
rect 65 14195 235 14365
rect 3085 1595 3255 1765
rect 3085 1955 3255 2125
rect 3085 2315 3255 2485
rect 3085 2675 3255 2845
rect 3085 3035 3255 3205
rect 3085 3395 3255 3565
rect 3085 3755 3255 3925
rect 3085 4115 3255 4285
rect 3085 4475 3255 4645
rect 3085 4835 3255 5005
rect 3085 5195 3255 5365
rect 3085 5555 3255 5725
rect 3085 5915 3255 6085
rect 3085 6275 3255 6445
rect 3085 6635 3255 6805
rect 3085 6995 3255 7165
rect 3085 7355 3255 7525
rect 425 515 595 685
rect 425 875 595 1045
rect 425 1235 595 1405
rect 425 1595 595 1765
rect 425 1955 595 2125
rect 425 2315 595 2485
rect 425 2675 595 2845
rect 425 3035 595 3205
rect 425 3395 595 3565
rect 425 3755 595 3925
rect 425 4115 595 4285
rect 425 4475 595 4645
rect 425 4835 595 5005
rect 425 5195 595 5365
rect 425 5555 595 5725
rect 425 5915 595 6085
rect 425 6275 595 6445
rect 425 6635 595 6805
rect 425 6995 595 7165
rect 425 7355 595 7525
rect 2725 2675 2895 2845
rect 2725 3035 2895 3205
rect 2725 3395 2895 3565
rect 2725 3755 2895 3925
rect 65 155 235 325
rect 65 515 235 685
rect 65 875 235 1045
rect 65 1235 235 1405
rect 65 1595 235 1765
rect 65 1955 235 2125
rect 65 2315 235 2485
rect 65 2675 235 2845
rect 65 3035 235 3205
rect 65 3395 235 3565
rect 65 3755 235 3925
rect 65 4115 235 4285
rect 65 4475 235 4645
rect 65 4835 235 5005
rect 65 5195 235 5365
rect 65 5555 235 5725
rect 65 5915 235 6085
rect 65 6275 235 6445
rect 65 6635 235 6805
rect 65 6995 235 7165
rect 65 7355 235 7525
rect 2725 4115 2895 4285
rect 2725 4475 2895 4645
rect 2725 4835 2895 5005
rect 2725 5195 2895 5365
rect 2725 5555 2895 5725
rect 2725 5915 2895 6085
rect 2725 6275 2895 6445
rect 2725 6635 2895 6805
rect 2725 6995 2895 7165
rect 2725 7355 2895 7525
rect 2725 1235 2895 1405
rect 2725 1595 2895 1765
rect 2725 1955 2895 2125
rect 2725 2315 2895 2485
rect 425 155 595 325
rect 3085 155 3255 325
rect 3085 515 3255 685
rect 3085 875 3255 1045
rect 3085 1235 3255 1405
rect 2725 155 2895 325
rect 2725 515 2895 685
rect 2725 875 2895 1045
<< l67d44 >>
rect 65 15275 235 15445
rect 425 15275 595 15445
rect 2725 15275 2895 15445
rect 3085 15275 3255 15445
rect 65 22835 235 23005
rect 425 22835 595 23005
rect 2725 22835 2895 23005
rect 3085 22835 3255 23005
rect 65 24275 235 24445
rect 65 24635 235 24805
rect 65 24995 235 25165
rect 65 25355 235 25525
rect 65 25715 235 25885
rect 65 26075 235 26245
rect 65 26435 235 26605
rect 65 26795 235 26965
rect 65 27155 235 27325
rect 65 27515 235 27685
rect 65 27875 235 28045
rect 65 28235 235 28405
rect 65 28595 235 28765
rect 65 28955 235 29125
rect 65 29315 235 29485
rect 65 29675 235 29845
rect 65 23195 235 23365
rect 425 23195 595 23365
rect 425 23555 595 23725
rect 425 23915 595 24085
rect 425 24275 595 24445
rect 425 24635 595 24805
rect 425 24995 595 25165
rect 425 25355 595 25525
rect 425 25715 595 25885
rect 425 26075 595 26245
rect 425 26435 595 26605
rect 425 26795 595 26965
rect 425 27155 595 27325
rect 425 27515 595 27685
rect 425 27875 595 28045
rect 425 28235 595 28405
rect 425 28595 595 28765
rect 425 28955 595 29125
rect 425 29315 595 29485
rect 425 29675 595 29845
rect 65 23555 235 23725
rect 2725 23195 2895 23365
rect 2725 23555 2895 23725
rect 2725 23915 2895 24085
rect 2725 24275 2895 24445
rect 2725 24635 2895 24805
rect 2725 24995 2895 25165
rect 2725 25355 2895 25525
rect 2725 25715 2895 25885
rect 2725 26075 2895 26245
rect 2725 26435 2895 26605
rect 2725 26795 2895 26965
rect 2725 27155 2895 27325
rect 2725 27515 2895 27685
rect 2725 27875 2895 28045
rect 2725 28235 2895 28405
rect 2725 28595 2895 28765
rect 2725 28955 2895 29125
rect 2725 29315 2895 29485
rect 2725 29675 2895 29845
rect 65 23915 235 24085
rect 3085 23195 3255 23365
rect 3085 23555 3255 23725
rect 3085 23915 3255 24085
rect 3085 24275 3255 24445
rect 3085 24635 3255 24805
rect 3085 24995 3255 25165
rect 3085 25355 3255 25525
rect 3085 25715 3255 25885
rect 3085 26075 3255 26245
rect 3085 26435 3255 26605
rect 3085 26795 3255 26965
rect 3085 27155 3255 27325
rect 3085 27515 3255 27685
rect 3085 27875 3255 28045
rect 3085 28235 3255 28405
rect 3085 28595 3255 28765
rect 3085 28955 3255 29125
rect 3085 29315 3255 29485
rect 3085 29675 3255 29845
rect 855 30280 1025 30450
rect 1215 30280 1385 30450
rect 1575 30280 1745 30450
rect 1935 30280 2105 30450
rect 2295 30280 2465 30450
rect 2725 17795 2895 17965
rect 2725 18155 2895 18325
rect 2725 18515 2895 18685
rect 2725 18875 2895 19045
rect 2725 19235 2895 19405
rect 2725 19595 2895 19765
rect 2725 19955 2895 20125
rect 2725 20315 2895 20485
rect 2725 20675 2895 20845
rect 2725 21035 2895 21205
rect 2725 21395 2895 21565
rect 2725 21755 2895 21925
rect 2725 22115 2895 22285
rect 2725 22475 2895 22645
rect 425 16355 595 16525
rect 425 16715 595 16885
rect 425 17075 595 17245
rect 425 17435 595 17605
rect 425 17795 595 17965
rect 425 18155 595 18325
rect 425 18515 595 18685
rect 425 18875 595 19045
rect 425 19235 595 19405
rect 425 19595 595 19765
rect 425 19955 595 20125
rect 425 20315 595 20485
rect 425 20675 595 20845
rect 425 21035 595 21205
rect 425 21395 595 21565
rect 425 21755 595 21925
rect 425 22115 595 22285
rect 425 22475 595 22645
rect 65 17795 235 17965
rect 65 18155 235 18325
rect 65 16355 235 16525
rect 3085 15635 3255 15805
rect 3085 15995 3255 16165
rect 3085 16355 3255 16525
rect 3085 16715 3255 16885
rect 3085 17075 3255 17245
rect 3085 17435 3255 17605
rect 3085 17795 3255 17965
rect 3085 18155 3255 18325
rect 3085 18515 3255 18685
rect 3085 18875 3255 19045
rect 3085 19235 3255 19405
rect 3085 19595 3255 19765
rect 3085 19955 3255 20125
rect 3085 20315 3255 20485
rect 3085 20675 3255 20845
rect 3085 21035 3255 21205
rect 3085 21395 3255 21565
rect 3085 21755 3255 21925
rect 3085 22115 3255 22285
rect 3085 22475 3255 22645
rect 65 18515 235 18685
rect 65 18875 235 19045
rect 65 19235 235 19405
rect 65 19595 235 19765
rect 65 19955 235 20125
rect 65 20315 235 20485
rect 65 20675 235 20845
rect 65 21035 235 21205
rect 65 21395 235 21565
rect 65 21755 235 21925
rect 65 22115 235 22285
rect 65 22475 235 22645
rect 65 16715 235 16885
rect 65 17075 235 17245
rect 65 17435 235 17605
rect 65 15635 235 15805
rect 425 15635 595 15805
rect 425 15995 595 16165
rect 65 15995 235 16165
rect 2725 15635 2895 15805
rect 2725 15995 2895 16165
rect 2725 16355 2895 16525
rect 2725 16715 2895 16885
rect 2725 17075 2895 17245
rect 2725 17435 2895 17605
rect 2725 7715 2895 7885
rect 425 7715 595 7885
rect 3085 7715 3255 7885
rect 65 7715 235 7885
rect 2725 9155 2895 9325
rect 2725 9515 2895 9685
rect 2725 9875 2895 10045
rect 2725 10235 2895 10405
rect 2725 10595 2895 10765
rect 2725 10955 2895 11125
rect 2725 11315 2895 11485
rect 2725 11675 2895 11845
rect 2725 12035 2895 12205
rect 2725 12395 2895 12565
rect 2725 12755 2895 12925
rect 2725 13115 2895 13285
rect 2725 13475 2895 13645
rect 2725 13835 2895 14005
rect 2725 14195 2895 14365
rect 2725 14555 2895 14725
rect 2725 14915 2895 15085
rect 65 14555 235 14725
rect 2725 8075 2895 8245
rect 425 8075 595 8245
rect 425 8435 595 8605
rect 425 8795 595 8965
rect 425 9155 595 9325
rect 425 9515 595 9685
rect 425 9875 595 10045
rect 425 10235 595 10405
rect 425 10595 595 10765
rect 425 10955 595 11125
rect 425 11315 595 11485
rect 425 11675 595 11845
rect 425 12035 595 12205
rect 425 12395 595 12565
rect 425 12755 595 12925
rect 425 13115 595 13285
rect 425 13475 595 13645
rect 425 13835 595 14005
rect 425 14195 595 14365
rect 2725 8435 2895 8605
rect 3085 8075 3255 8245
rect 3085 8435 3255 8605
rect 3085 8795 3255 8965
rect 3085 9155 3255 9325
rect 3085 9515 3255 9685
rect 3085 9875 3255 10045
rect 3085 10235 3255 10405
rect 3085 10595 3255 10765
rect 3085 10955 3255 11125
rect 3085 11315 3255 11485
rect 3085 11675 3255 11845
rect 3085 12035 3255 12205
rect 3085 12395 3255 12565
rect 3085 12755 3255 12925
rect 3085 13115 3255 13285
rect 3085 13475 3255 13645
rect 3085 13835 3255 14005
rect 3085 14195 3255 14365
rect 3085 14555 3255 14725
rect 3085 14915 3255 15085
rect 425 14555 595 14725
rect 425 14915 595 15085
rect 65 14915 235 15085
rect 2725 8795 2895 8965
rect 65 8075 235 8245
rect 65 8435 235 8605
rect 65 8795 235 8965
rect 65 9155 235 9325
rect 65 9515 235 9685
rect 65 9875 235 10045
rect 65 10235 235 10405
rect 65 10595 235 10765
rect 65 10955 235 11125
rect 65 11315 235 11485
rect 65 11675 235 11845
rect 65 12035 235 12205
rect 65 12395 235 12565
rect 65 12755 235 12925
rect 65 13115 235 13285
rect 65 13475 235 13645
rect 65 13835 235 14005
rect 65 14195 235 14365
rect 3085 1595 3255 1765
rect 3085 1955 3255 2125
rect 3085 2315 3255 2485
rect 3085 2675 3255 2845
rect 3085 3035 3255 3205
rect 3085 3395 3255 3565
rect 3085 3755 3255 3925
rect 3085 4115 3255 4285
rect 3085 4475 3255 4645
rect 3085 4835 3255 5005
rect 3085 5195 3255 5365
rect 3085 5555 3255 5725
rect 3085 5915 3255 6085
rect 3085 6275 3255 6445
rect 3085 6635 3255 6805
rect 3085 6995 3255 7165
rect 3085 7355 3255 7525
rect 425 515 595 685
rect 425 875 595 1045
rect 425 1235 595 1405
rect 425 1595 595 1765
rect 425 1955 595 2125
rect 425 2315 595 2485
rect 425 2675 595 2845
rect 425 3035 595 3205
rect 425 3395 595 3565
rect 425 3755 595 3925
rect 425 4115 595 4285
rect 425 4475 595 4645
rect 425 4835 595 5005
rect 425 5195 595 5365
rect 425 5555 595 5725
rect 425 5915 595 6085
rect 425 6275 595 6445
rect 425 6635 595 6805
rect 425 6995 595 7165
rect 425 7355 595 7525
rect 2725 2675 2895 2845
rect 2725 3035 2895 3205
rect 2725 3395 2895 3565
rect 2725 3755 2895 3925
rect 65 155 235 325
rect 65 515 235 685
rect 65 875 235 1045
rect 65 1235 235 1405
rect 65 1595 235 1765
rect 65 1955 235 2125
rect 65 2315 235 2485
rect 65 2675 235 2845
rect 65 3035 235 3205
rect 65 3395 235 3565
rect 65 3755 235 3925
rect 65 4115 235 4285
rect 65 4475 235 4645
rect 65 4835 235 5005
rect 65 5195 235 5365
rect 65 5555 235 5725
rect 65 5915 235 6085
rect 65 6275 235 6445
rect 65 6635 235 6805
rect 65 6995 235 7165
rect 65 7355 235 7525
rect 2725 4115 2895 4285
rect 2725 4475 2895 4645
rect 2725 4835 2895 5005
rect 2725 5195 2895 5365
rect 2725 5555 2895 5725
rect 2725 5915 2895 6085
rect 2725 6275 2895 6445
rect 2725 6635 2895 6805
rect 2725 6995 2895 7165
rect 2725 7355 2895 7525
rect 2725 1235 2895 1405
rect 2725 1595 2895 1765
rect 2725 1955 2895 2125
rect 2725 2315 2895 2485
rect 425 155 595 325
rect 3085 155 3255 325
rect 3085 515 3255 685
rect 3085 875 3255 1045
rect 3085 1235 3255 1405
rect 2725 155 2895 325
rect 2725 515 2895 685
rect 2725 875 2895 1045
<< l95d20 >>
rect 650 30190 2670 30540
<< l67d20 >>
rect 65 75 595 29925
rect 2725 75 3255 29925
rect 775 30280 2545 30450
<< l68d20 >>
rect 35 95 625 29905
rect 2695 95 3285 29905
rect 795 30250 2525 30480
<< l65d20 >>
rect 0 0 3320 30000
<< l93d44 >>
rect -125 -125 3445 30125
<< end >>
