magic
tech sky130A
magscale 1 2
timestamp 1698900908
<< error_s >>
rect 17140 21212 17152 21218
rect 17163 21194 17164 21206
rect 20416 21122 20422 21128
rect 20386 21098 20392 21118
rect 20344 21010 20350 21030
rect 20386 20988 20392 20994
rect 17163 20826 17164 20838
rect 17140 20814 17152 20820
rect 21874 20722 21875 20900
rect 21915 20722 21916 20900
rect 21874 20538 21875 20652
rect 21804 20469 21875 20538
rect 21915 20538 21916 20652
rect 21915 20469 21986 20538
rect 21915 20468 21917 20469
rect 21916 20467 21944 20468
rect 2298 20388 2498 20410
rect 21874 20398 21875 20467
rect 21915 20398 21944 20467
rect 21915 20397 21917 20398
rect 11340 20008 11540 20030
rect 21874 19966 21875 20397
rect 21915 19966 21916 20397
rect 22371 20284 22372 20646
rect 22301 20215 22372 20284
rect 22412 20284 22413 20646
rect 22868 20538 22869 20900
rect 22798 20469 22869 20538
rect 22909 20538 22910 20900
rect 22909 20469 22980 20538
rect 22909 20468 22911 20469
rect 22910 20467 22938 20468
rect 22868 20398 22869 20467
rect 22909 20398 22938 20467
rect 22909 20397 22911 20398
rect 22412 20215 22483 20284
rect 22412 20214 22414 20215
rect 22413 20213 22441 20214
rect 22371 20144 22372 20213
rect 22412 20144 22441 20213
rect 22412 20143 22414 20144
rect 22371 19712 22372 20143
rect 22412 19712 22413 20143
rect 22868 19966 22869 20397
rect 22909 19966 22910 20397
rect 23365 20284 23366 20646
rect 23295 20215 23366 20284
rect 23406 20284 23407 20646
rect 23862 20538 23863 20900
rect 23792 20469 23863 20538
rect 23903 20538 23904 20900
rect 23903 20469 23974 20538
rect 23903 20468 23905 20469
rect 23904 20467 23932 20468
rect 23862 20398 23863 20467
rect 23903 20398 23932 20467
rect 23903 20397 23905 20398
rect 23406 20215 23477 20284
rect 23406 20214 23408 20215
rect 23407 20213 23435 20214
rect 23365 20144 23366 20213
rect 23406 20144 23435 20213
rect 23406 20143 23408 20144
rect 23365 19712 23366 20143
rect 23406 19712 23407 20143
rect 23862 19966 23863 20397
rect 23903 19966 23904 20397
rect 24359 20284 24360 20646
rect 24289 20215 24360 20284
rect 24400 20284 24401 20646
rect 24856 20538 24857 20900
rect 24786 20469 24857 20538
rect 24897 20538 24898 20900
rect 24897 20469 24968 20538
rect 24897 20468 24899 20469
rect 24898 20467 24926 20468
rect 24856 20398 24857 20467
rect 24897 20398 24926 20467
rect 24897 20397 24899 20398
rect 24400 20215 24471 20284
rect 24400 20214 24402 20215
rect 24401 20213 24429 20214
rect 24359 20144 24360 20213
rect 24400 20144 24429 20213
rect 24400 20143 24402 20144
rect 24359 19712 24360 20143
rect 24400 19712 24401 20143
rect 24856 19966 24857 20397
rect 24897 19966 24898 20397
rect 25353 20284 25354 20646
rect 25283 20215 25354 20284
rect 25394 20284 25395 20646
rect 25394 20215 25465 20284
rect 25394 20214 25396 20215
rect 25395 20213 25423 20214
rect 25353 20144 25354 20213
rect 25394 20144 25423 20213
rect 25394 20143 25396 20144
rect 25353 19712 25354 20143
rect 25394 19712 25395 20143
rect 2288 19666 8340 19667
rect 11330 19286 17382 19287
rect 21302 17852 21345 17920
rect 1317 9586 1339 9824
rect 2006 9586 2049 15654
rect 21344 11826 21345 17852
rect 22066 17668 22088 17868
rect 2006 9560 2007 9586
rect 2527 1366 2549 1604
rect 3216 1366 3259 7434
rect 14969 4073 21105 4116
rect 4668 3749 4811 4003
rect 4922 2154 5065 3749
rect 20799 3384 21037 3406
rect 6930 2154 13066 2197
rect 12760 1465 12998 1487
rect 3216 1340 3217 1366
<< metal1 >>
rect 1856 20837 11335 21273
rect 400 20400 2293 20837
rect 400 9565 836 20400
rect 1856 17575 2264 20197
rect 10898 20020 11335 20837
rect 16983 21212 17057 21786
rect 21755 21726 22025 21786
rect 22252 21726 22577 21786
rect 22749 21726 23129 21786
rect 23246 21726 23681 21786
rect 24159 21726 24520 21786
rect 24711 21726 25017 21786
rect 25263 21726 25514 21786
rect 25815 21726 26011 21786
rect 16983 20820 17108 21212
rect 20526 21017 20645 21091
rect 10303 19409 11191 19817
rect 20571 19437 20645 21017
rect 21755 20772 21815 21726
rect 22252 21026 22312 21726
rect 22749 21280 22809 21726
rect 23246 21534 23306 21726
rect 22885 21474 23306 21534
rect 24460 21534 24520 21726
rect 24460 21474 24881 21534
rect 22388 21220 22809 21280
rect 24957 21280 25017 21726
rect 24957 21220 25378 21280
rect 21891 20966 22312 21026
rect 25454 21026 25514 21726
rect 25454 20966 25875 21026
rect 21394 20712 21815 20772
rect 25951 20772 26011 21726
rect 25951 20712 26372 20772
rect 19345 19029 20645 19437
rect 20291 18017 20571 19029
rect 21925 18310 22362 20154
rect 21925 17873 22964 18310
rect 400 9128 1273 9565
rect 1476 9128 3474 9536
rect 836 1345 1273 9128
rect 836 908 2483 1345
rect 5009 1316 5417 2004
rect 13048 1624 13456 3923
rect 21087 3543 21495 9863
rect 22527 3339 22964 17873
rect 21058 2903 22964 3339
rect 21058 1421 21495 2903
rect 2686 1016 5417 1316
rect 13019 984 21495 1421
rect 13019 908 13456 984
rect 2046 472 13456 908
<< metal2 >>
rect 0 21370 3864 22304
rect 27916 22260 31464 22304
rect 8702 21370 16506 22085
rect 27916 21370 31116 22260
rect 0 21116 31116 21370
rect 0 20290 16692 21116
rect 20897 20828 31116 21116
rect 20897 20290 21026 20828
rect 21437 20461 21871 20470
rect 21437 20405 21446 20461
rect 21502 20405 21536 20461
rect 21592 20405 21626 20461
rect 21682 20405 21716 20461
rect 21772 20405 21806 20461
rect 21862 20405 21871 20461
rect 21437 20396 21871 20405
rect 0 20005 21026 20290
rect 22225 20005 31116 20828
rect 0 18754 31116 20005
rect 0 17854 1919 18754
rect 10697 18393 31116 18754
rect 0 9252 2904 17854
rect 10697 17755 10970 18393
rect 3909 17367 10970 17755
rect 3909 9770 19400 17367
rect 3909 9252 4122 9770
rect 5132 9461 19400 9770
rect 20449 9461 31116 18393
rect 0 1079 4122 9252
rect 5132 5988 31116 9461
rect 5132 4955 12636 5988
rect 21449 4955 31116 5988
rect 5132 4086 31116 4955
rect 13400 3056 31116 4086
rect 5132 1079 31116 3056
rect 0 44 31116 1079
rect 31412 44 31464 22260
rect 0 0 31464 44
<< via2 >>
rect 17125 20716 17181 20772
rect 17205 20716 17261 20772
rect 17285 20716 17341 20772
rect 17365 20716 17421 20772
rect 17445 20716 17501 20772
rect 17525 20716 17581 20772
rect 17605 20716 17661 20772
rect 17685 20716 17741 20772
rect 17765 20716 17821 20772
rect 17845 20716 17901 20772
rect 17925 20716 17981 20772
rect 18005 20716 18061 20772
rect 18085 20716 18141 20772
rect 18165 20716 18221 20772
rect 18245 20716 18301 20772
rect 18325 20716 18381 20772
rect 18405 20716 18461 20772
rect 18485 20716 18541 20772
rect 18565 20716 18621 20772
rect 18645 20716 18701 20772
rect 18725 20716 18781 20772
rect 18805 20716 18861 20772
rect 18885 20716 18941 20772
rect 18965 20716 19021 20772
rect 19045 20716 19101 20772
rect 19125 20716 19181 20772
rect 19205 20716 19261 20772
rect 19285 20716 19341 20772
rect 19365 20716 19421 20772
rect 19445 20716 19501 20772
rect 19525 20716 19581 20772
rect 19605 20716 19661 20772
rect 19685 20716 19741 20772
rect 19765 20716 19821 20772
rect 19845 20716 19901 20772
rect 19925 20716 19981 20772
rect 20005 20716 20061 20772
rect 20085 20716 20141 20772
rect 20165 20716 20221 20772
rect 20245 20716 20301 20772
rect 20325 20716 20381 20772
rect 20405 20716 20461 20772
rect 21446 20405 21502 20461
rect 21536 20405 21592 20461
rect 21626 20405 21682 20461
rect 21716 20405 21772 20461
rect 21806 20405 21862 20461
rect 2366 18197 10262 18333
rect 11408 17817 19304 17953
rect 3340 9638 3476 17534
rect 19875 9904 20011 17800
rect 4550 1418 4686 9314
rect 13089 5406 20985 5542
rect 5050 3488 12946 3624
rect 31116 44 31412 22260
<< metal3 >>
rect 0 22264 8226 22304
rect 0 40 48 22264
rect 352 21370 8226 22264
rect 27916 21370 30633 22304
rect 352 20772 30633 21370
rect 352 20716 17125 20772
rect 17181 20716 17205 20772
rect 17261 20716 17285 20772
rect 17341 20716 17365 20772
rect 17421 20716 17445 20772
rect 17501 20716 17525 20772
rect 17581 20716 17605 20772
rect 17661 20716 17685 20772
rect 17741 20716 17765 20772
rect 17821 20716 17845 20772
rect 17901 20716 17925 20772
rect 17981 20716 18005 20772
rect 18061 20716 18085 20772
rect 18141 20716 18165 20772
rect 18221 20716 18245 20772
rect 18301 20716 18325 20772
rect 18381 20716 18405 20772
rect 18461 20716 18485 20772
rect 18541 20716 18565 20772
rect 18621 20716 18645 20772
rect 18701 20716 18725 20772
rect 18781 20716 18805 20772
rect 18861 20716 18885 20772
rect 18941 20716 18965 20772
rect 19021 20716 19045 20772
rect 19101 20716 19125 20772
rect 19181 20716 19205 20772
rect 19261 20716 19285 20772
rect 19341 20716 19365 20772
rect 19421 20716 19445 20772
rect 19501 20716 19525 20772
rect 19581 20716 19605 20772
rect 19661 20716 19685 20772
rect 19741 20716 19765 20772
rect 19821 20716 19845 20772
rect 19901 20716 19925 20772
rect 19981 20716 20005 20772
rect 20061 20716 20085 20772
rect 20141 20716 20165 20772
rect 20221 20716 20245 20772
rect 20301 20716 20325 20772
rect 20381 20716 20405 20772
rect 20461 20716 30633 20772
rect 352 20461 30633 20716
rect 352 20405 21446 20461
rect 21502 20405 21536 20461
rect 21592 20405 21626 20461
rect 21682 20405 21716 20461
rect 21772 20405 21806 20461
rect 21862 20405 30633 20461
rect 352 18333 30633 20405
rect 352 18197 2366 18333
rect 10262 18197 30633 18333
rect 352 17953 30633 18197
rect 352 17817 11408 17953
rect 19304 17817 30633 17953
rect 352 17800 30633 17817
rect 352 17534 19875 17800
rect 352 9638 3340 17534
rect 3476 9904 19875 17534
rect 20011 9904 30633 17800
rect 3476 9638 30633 9904
rect 352 9314 30633 9638
rect 352 1418 4550 9314
rect 4686 5542 30633 9314
rect 4686 5406 13089 5542
rect 20985 5406 30633 5542
rect 4686 3624 30633 5406
rect 4686 3488 5050 3624
rect 12946 3488 30633 3624
rect 4686 1418 30633 3488
rect 352 40 30633 1418
rect 0 0 30633 40
rect 31064 22264 31464 22304
rect 31064 40 31112 22264
rect 31416 40 31464 22264
rect 31064 0 31464 40
<< via3 >>
rect 48 40 352 22264
rect 31112 22260 31416 22264
rect 31112 44 31116 22260
rect 31116 44 31412 22260
rect 31412 44 31416 22260
rect 31112 40 31416 44
<< metal4 >>
rect 0 22264 400 22304
rect 0 40 48 22264
rect 352 40 400 22264
rect 4294 22104 4354 22304
rect 4846 22104 4906 22304
rect 5398 22104 5458 22304
rect 5950 22104 6010 22304
rect 6502 22104 6562 22304
rect 7054 22104 7114 22304
rect 7606 22104 7666 22304
rect 8158 22104 8218 22304
rect 8710 22104 8770 22304
rect 9262 22104 9322 22304
rect 9814 22104 9874 22304
rect 10366 22104 10426 22304
rect 10918 22104 10978 22304
rect 11470 22104 11530 22304
rect 12022 22104 12082 22304
rect 12574 22104 12634 22304
rect 13126 22104 13186 22304
rect 13678 22104 13738 22304
rect 14230 22104 14290 22304
rect 14782 22104 14842 22304
rect 15334 22104 15394 22304
rect 15886 22104 15946 22304
rect 16438 22104 16498 22304
rect 16990 22104 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22104 22018 22304
rect 22510 22104 22570 22304
rect 23062 22104 23122 22304
rect 23614 22104 23674 22304
rect 24166 22104 24226 22304
rect 24718 22104 24778 22304
rect 25270 22104 25330 22304
rect 25822 22104 25882 22304
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 31064 22264 31464 22304
rect 0 0 400 40
rect 31064 40 31112 22264
rect 31416 40 31464 22264
rect 31064 0 31464 40
use dac_8bit  dac_8bit_0
timestamp 1698900908
transform 0 -1 26400 -1 0 21506
box 22 22 1794 5012
use driver  driver_0
timestamp 1698900908
transform -1 0 61693 0 -1 61377
box 41155 40041 44640 40681
use inv_strvd  inv_strvd_0
timestamp 1698900908
transform 0 1 2378 1 0 5319
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_1
timestamp 1698900908
transform 1 0 6267 0 -1 20505
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_2
timestamp 1698900908
transform 1 0 15309 0 -1 20125
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_3
timestamp 1698900908
transform -1 0 9045 0 1 1316
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_4
timestamp 1698900908
transform 0 -1 22183 -1 0 13899
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_5
timestamp 1698900908
transform 0 1 1168 1 0 13539
box -4118 -159 4123 2433
use inv_strvd  inv_strvd_6
timestamp 1698900908
transform -1 0 17084 0 1 3235
box -4118 -159 4123 2433
use pin_connect  pin_connect_0
timestamp 1698900908
transform 1 0 27471 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_1
timestamp 1698900908
transform 1 0 26919 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_2
timestamp 1698900908
transform 1 0 26367 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_3
timestamp 1698900908
transform 1 0 25815 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_4
timestamp 1698900908
transform 1 0 25263 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_5
timestamp 1698900908
transform 1 0 24711 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_6
timestamp 1698900908
transform 1 0 24159 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_7
timestamp 1698900908
transform 1 0 23607 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_8
timestamp 1698900908
transform 1 0 23055 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_9
timestamp 1698900908
transform 1 0 22503 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_10
timestamp 1698900908
transform 1 0 21951 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_11
timestamp 1698900908
transform 1 0 21399 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_12
timestamp 1698900908
transform 1 0 20847 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_13
timestamp 1698900908
transform 1 0 20295 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_14
timestamp 1698900908
transform 1 0 19743 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_15
timestamp 1698900908
transform 1 0 19191 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_16
timestamp 1698900908
transform 1 0 18639 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_17
timestamp 1698900908
transform 1 0 18087 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_18
timestamp 1698900908
transform 1 0 17535 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_19
timestamp 1698900908
transform 1 0 16983 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_20
timestamp 1698900908
transform 1 0 16431 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_21
timestamp 1698900908
transform 1 0 15879 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_22
timestamp 1698900908
transform 1 0 15327 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_23
timestamp 1698900908
transform 1 0 14775 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_24
timestamp 1698900908
transform 1 0 14223 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_25
timestamp 1698900908
transform 1 0 13671 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_26
timestamp 1698900908
transform 1 0 13119 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_27
timestamp 1698900908
transform 1 0 12567 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_28
timestamp 1698900908
transform 1 0 12015 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_29
timestamp 1698900908
transform 1 0 11463 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_30
timestamp 1698900908
transform 1 0 10911 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_31
timestamp 1698900908
transform 1 0 10359 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_32
timestamp 1698900908
transform 1 0 9807 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_33
timestamp 1698900908
transform 1 0 9255 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_34
timestamp 1698900908
transform 1 0 8703 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_35
timestamp 1698900908
transform 1 0 8151 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_36
timestamp 1698900908
transform 1 0 7599 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_37
timestamp 1698900908
transform 1 0 7047 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_38
timestamp 1698900908
transform 1 0 6495 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_39
timestamp 1698900908
transform 1 0 5943 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_40
timestamp 1698900908
transform 1 0 5391 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_41
timestamp 1698900908
transform 1 0 4839 0 1 21786
box -1 0 75 518
use pin_connect  pin_connect_42
timestamp 1698900908
transform 1 0 4287 0 1 21786
box -1 0 75 518
use tt_um_template  tt_um_template_0
timestamp 1698900908
transform 1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel metal4 s 31064 0 31464 22304 0 FreeSans 2000 0 0 0 VGND
port 2 nsew
rlabel metal4 s 26926 22104 26986 22304 4 clk
port 3 nsew
rlabel metal4 s 27478 22104 27538 22304 4 ena
port 4 nsew
rlabel metal4 s 26374 22104 26434 22304 4 rst_n
port 5 nsew
rlabel metal4 s 25822 22104 25882 22304 4 ui_in[0]
port 6 nsew
rlabel metal4 s 25270 22104 25330 22304 4 ui_in[1]
port 7 nsew
rlabel metal4 s 24718 22104 24778 22304 4 ui_in[2]
port 8 nsew
rlabel metal4 s 24166 22104 24226 22304 4 ui_in[3]
port 9 nsew
rlabel metal4 s 23614 22104 23674 22304 4 ui_in[4]
port 10 nsew
rlabel metal4 s 23062 22104 23122 22304 4 ui_in[5]
port 11 nsew
rlabel metal4 s 22510 22104 22570 22304 4 ui_in[6]
port 12 nsew
rlabel metal4 s 21958 22104 22018 22304 4 ui_in[7]
port 13 nsew
rlabel metal4 s 21406 22104 21466 22304 4 uio_in[0]
port 14 nsew
rlabel metal4 s 20854 22104 20914 22304 4 uio_in[1]
port 15 nsew
rlabel metal4 s 20302 22104 20362 22304 4 uio_in[2]
port 16 nsew
rlabel metal4 s 19750 22104 19810 22304 4 uio_in[3]
port 17 nsew
rlabel metal4 s 19198 22104 19258 22304 4 uio_in[4]
port 18 nsew
rlabel metal4 s 18646 22104 18706 22304 4 uio_in[5]
port 19 nsew
rlabel metal4 s 18094 22104 18154 22304 4 uio_in[6]
port 20 nsew
rlabel metal4 s 17542 22104 17602 22304 4 uio_in[7]
port 21 nsew
rlabel metal4 s 8158 22104 8218 22304 4 uio_oe[0]
port 22 nsew
rlabel metal4 s 7606 22104 7666 22304 4 uio_oe[1]
port 23 nsew
rlabel metal4 s 7054 22104 7114 22304 4 uio_oe[2]
port 24 nsew
rlabel metal4 s 6502 22104 6562 22304 4 uio_oe[3]
port 25 nsew
rlabel metal4 s 5950 22104 6010 22304 4 uio_oe[4]
port 26 nsew
rlabel metal4 s 5398 22104 5458 22304 4 uio_oe[5]
port 27 nsew
rlabel metal4 s 4846 22104 4906 22304 4 uio_oe[6]
port 28 nsew
rlabel metal4 s 4294 22104 4354 22304 4 uio_oe[7]
port 29 nsew
rlabel metal4 s 12574 22104 12634 22304 4 uio_out[0]
port 30 nsew
rlabel metal4 s 12022 22104 12082 22304 4 uio_out[1]
port 31 nsew
rlabel metal4 s 11470 22104 11530 22304 4 uio_out[2]
port 32 nsew
rlabel metal4 s 10918 22104 10978 22304 4 uio_out[3]
port 33 nsew
rlabel metal4 s 10366 22104 10426 22304 4 uio_out[4]
port 34 nsew
rlabel metal4 s 9814 22104 9874 22304 4 uio_out[5]
port 35 nsew
rlabel metal4 s 9262 22104 9322 22304 4 uio_out[6]
port 36 nsew
rlabel metal4 s 8710 22104 8770 22304 4 uio_out[7]
port 37 nsew
rlabel metal4 s 16990 22104 17050 22304 4 uo_out[0]
port 38 nsew
rlabel metal4 s 16438 22104 16498 22304 4 uo_out[1]
port 39 nsew
rlabel metal4 s 15886 22104 15946 22304 4 uo_out[2]
port 40 nsew
rlabel metal4 s 15334 22104 15394 22304 4 uo_out[3]
port 41 nsew
rlabel metal4 s 14782 22104 14842 22304 4 uo_out[4]
port 42 nsew
rlabel metal4 s 14230 22104 14290 22304 4 uo_out[5]
port 43 nsew
rlabel metal4 s 13678 22104 13738 22304 4 uo_out[6]
port 44 nsew
rlabel metal4 s 13126 22104 13186 22304 4 uo_out[7]
port 45 nsew
flabel metal4 s 0 0 400 22304 0 FreeSans 2000 0 0 0 VPWR
port 46 nsew
<< end >>
