magic
tech sky130a
timestamp 1698899266
<< checkpaint >>
rect 0 0 157320 111520
<< l68d20 >>
rect 112637 14515 114819 89365
rect 65096 4921 105291 7104
rect 1998 47823 4181 104185
rect 102854 95145 103224 105087
rect 111260 108628 112885 108928
rect 11464 104185 56674 106367
rect 109456 104832 111560 105132
rect 111941 106102 114045 106402
rect 108775 108628 110125 108928
rect 113745 108628 115645 108928
rect 126315 108628 127572 108928
rect 123555 108628 125087 108928
rect 114426 107372 116530 107672
rect 116230 108628 118405 108928
rect 127272 104832 129376 105132
rect 129757 103562 131861 103862
rect 129075 108628 130057 108928
rect 120795 108628 122602 108928
rect 129757 103862 130057 108628
rect 124787 106402 125087 108628
rect 122302 107372 124406 107672
rect 127272 105132 127572 108628
rect 124787 106102 126891 106402
rect 122302 107672 122602 108628
rect 116230 107672 116530 108628
rect 113745 106402 114045 108628
rect 111260 105132 111560 108628
rect 108775 103862 109075 108628
rect 106971 103562 109075 103862
rect 102628 105087 103224 105457
rect 84915 104102 85285 108928
rect 85285 104102 85542 106062
rect 96725 95145 102854 97185
rect 101453 90084 102854 95145
rect 111810 89365 114819 91548
rect 109627 89365 111810 100772
rect 51515 97045 55955 99085
rect 4181 102002 11464 104185
rect 9282 104185 11464 106367
rect 54491 100102 56674 104185
rect 9280 87874 11320 100985
rect 13430 5079 27085 6579
rect 65240 8121 67280 19614
rect 12413 2358 65096 4541
rect 10230 2358 12413 4541
rect 4181 4541 12413 6723
rect 4181 6723 6363 47823
rect 1998 45640 4181 47823
rect 65096 2358 67278 4921
rect 7380 45639 17370 47679
rect 25045 6579 27085 10021
rect 105291 14515 112637 16697
rect 105291 4921 107474 14515
rect 105435 17714 107475 49314
<< l69d20 >>
rect 67000 0 107243 24776
rect 0 0 14522 89271
rect 19322 93769 54851 106848
rect 21507 48852 96998 86834
rect 63180 29938 96998 48852
rect 43510 106848 82530 110423
rect 0 93769 19322 111520
rect 14522 5395 20612 46258
rect 83462 91965 105129 101449
rect 104483 101449 105129 104142
rect 96998 29938 107243 47306
rect 102245 47306 107243 91965
rect 0 89271 9593 93769
rect 19544 86834 53483 88775
rect 19544 48852 21507 86834
rect 19544 46258 20612 48852
rect 53483 86834 54851 93769
rect 63180 20430 67000 24776
rect 105129 91965 107243 100027
rect 14522 0 25661 5395
rect 139578 100027 157320 111520
rect 107186 101982 109356 102352
rect 25661 0 67000 15279
rect 25661 20430 63180 48852
rect 111126 100027 139578 104142
rect 104483 104142 139578 106848
rect 107243 0 157320 100027
rect 54851 91965 83462 106848
rect 83462 105582 104483 106848
<< l70d44 >>
rect 155620 83460 155820 83660
rect 156820 83460 157020 83660
rect 156420 83460 156620 83660
rect 156020 83460 156220 83660
rect 155620 104260 155820 104460
rect 156420 104260 156620 104460
rect 156020 104260 156220 104460
rect 156820 104260 157020 104460
rect 156820 107860 157020 108060
rect 156020 110660 156220 110860
rect 156820 108260 157020 108460
rect 156020 111060 156220 111260
rect 156820 108660 157020 108860
rect 156820 109060 157020 109260
rect 156820 109460 157020 109660
rect 156820 109860 157020 110060
rect 156820 110260 157020 110460
rect 156020 108660 156220 108860
rect 156820 110660 157020 110860
rect 155620 104660 155820 104860
rect 156820 111060 157020 111260
rect 155620 105060 155820 105260
rect 155620 105460 155820 105660
rect 155620 105860 155820 106060
rect 155620 106260 155820 106460
rect 155620 106660 155820 106860
rect 156820 106260 157020 106460
rect 155620 107060 155820 107260
rect 156420 104660 156620 104860
rect 155620 107460 155820 107660
rect 156420 105060 156620 105260
rect 155620 107860 155820 108060
rect 156420 105460 156620 105660
rect 155620 108260 155820 108460
rect 156420 105860 156620 106060
rect 156020 109460 156220 109660
rect 155620 108660 155820 108860
rect 156420 106260 156620 106460
rect 155620 109060 155820 109260
rect 156420 106660 156620 106860
rect 155620 109460 155820 109660
rect 156420 107060 156620 107260
rect 155620 109860 155820 110060
rect 156420 107460 156620 107660
rect 155620 110260 155820 110460
rect 156420 107860 156620 108060
rect 155620 110660 155820 110860
rect 156420 108260 156620 108460
rect 155620 111060 155820 111260
rect 156420 108660 156620 108860
rect 156420 109060 156620 109260
rect 156420 109460 156620 109660
rect 156420 109860 156620 110060
rect 156420 110260 156620 110460
rect 156420 110660 156620 110860
rect 156420 111060 156620 111260
rect 156020 109060 156220 109260
rect 156020 104660 156220 104860
rect 156020 105060 156220 105260
rect 156020 105460 156220 105660
rect 156020 105860 156220 106060
rect 156020 106260 156220 106460
rect 156020 106660 156220 106860
rect 156820 106660 157020 106860
rect 156020 107060 156220 107260
rect 156820 104660 157020 104860
rect 156020 107460 156220 107660
rect 156820 105060 157020 105260
rect 156020 107860 156220 108060
rect 156820 105460 157020 105660
rect 156020 108260 156220 108460
rect 156820 105860 157020 106060
rect 156820 107060 157020 107260
rect 156020 109860 156220 110060
rect 156820 107460 157020 107660
rect 156020 110260 156220 110460
rect 156020 99060 156220 99260
rect 156420 98660 156620 98860
rect 156820 102660 157020 102860
rect 155620 101460 155820 101660
rect 156420 97460 156620 97660
rect 156420 99060 156620 99260
rect 156020 99460 156220 99660
rect 155620 101860 155820 102060
rect 156820 103060 157020 103260
rect 156420 99460 156620 99660
rect 155620 99860 155820 100060
rect 155620 102260 155820 102460
rect 156020 99860 156220 100060
rect 156420 99860 156620 100060
rect 155620 102660 155820 102860
rect 156820 103460 157020 103660
rect 156420 100260 156620 100460
rect 155620 103060 155820 103260
rect 156020 100260 156220 100460
rect 156420 100660 156620 100860
rect 155620 103460 155820 103660
rect 155620 98660 155820 98860
rect 156420 101060 156620 101260
rect 155620 103860 155820 104060
rect 156420 97860 156620 98060
rect 156020 100660 156220 100860
rect 156420 101460 156620 101660
rect 155620 97460 155820 97660
rect 156020 101060 156220 101260
rect 156420 101860 156620 102060
rect 156820 97460 157020 97660
rect 156820 103860 157020 104060
rect 156420 102260 156620 102460
rect 156820 97860 157020 98060
rect 156420 102660 156620 102860
rect 156020 101460 156220 101660
rect 156420 103060 156620 103260
rect 156820 98260 157020 98460
rect 156420 103460 156620 103660
rect 155620 99460 155820 99660
rect 156420 103860 156620 104060
rect 156020 101860 156220 102060
rect 156820 98660 157020 98860
rect 155620 97860 155820 98060
rect 156020 102260 156220 102460
rect 156820 99060 157020 99260
rect 156020 102660 156220 102860
rect 156820 99460 157020 99660
rect 156820 99860 157020 100060
rect 156020 103060 156220 103260
rect 156820 100260 157020 100460
rect 156020 103460 156220 103660
rect 156820 100660 157020 100860
rect 156020 103860 156220 104060
rect 156020 97460 156220 97660
rect 156820 101060 157020 101260
rect 155620 100660 155820 100860
rect 156020 97860 156220 98060
rect 155620 100260 155820 100460
rect 156820 101460 157020 101660
rect 156020 98260 156220 98460
rect 156820 101860 157020 102060
rect 155620 99060 155820 99260
rect 156020 98660 156220 98860
rect 156820 102260 157020 102460
rect 156420 98260 156620 98460
rect 155620 98260 155820 98460
rect 155620 101060 155820 101260
rect 155620 90260 155820 90460
rect 156020 90260 156220 90460
rect 156820 90260 157020 90460
rect 156420 90260 156620 90460
rect 155620 92660 155820 92860
rect 156020 94660 156220 94860
rect 155620 96260 155820 96460
rect 156020 95060 156220 95260
rect 156420 94660 156620 94860
rect 156420 95460 156620 95660
rect 156020 95460 156220 95660
rect 155620 93060 155820 93260
rect 156820 90660 157020 90860
rect 156420 93860 156620 94060
rect 156020 95860 156220 96060
rect 156820 91060 157020 91260
rect 156020 96260 156220 96460
rect 156820 91460 157020 91660
rect 155620 93460 155820 93660
rect 156820 91860 157020 92060
rect 156020 96660 156220 96860
rect 155620 96660 155820 96860
rect 156820 92260 157020 92460
rect 156420 91860 156620 92060
rect 156020 97060 156220 97260
rect 156420 94260 156620 94460
rect 156820 92660 157020 92860
rect 155620 93860 155820 94060
rect 156420 90660 156620 90860
rect 156820 93060 157020 93260
rect 156420 91060 156620 91260
rect 155620 94260 155820 94460
rect 156820 93460 157020 93660
rect 155620 97060 155820 97260
rect 156820 93860 157020 94060
rect 156420 91460 156620 91660
rect 156020 93860 156220 94060
rect 156420 93460 156620 93660
rect 156420 96260 156620 96460
rect 156020 94260 156220 94460
rect 156020 91060 156220 91260
rect 155620 95460 155820 95660
rect 155620 91060 155820 91260
rect 156020 91460 156220 91660
rect 156820 96260 157020 96460
rect 156420 92660 156620 92860
rect 156020 91860 156220 92060
rect 155620 91460 155820 91660
rect 156820 96660 157020 96860
rect 156020 92260 156220 92460
rect 156420 96660 156620 96860
rect 155620 91860 155820 92060
rect 156020 92660 156220 92860
rect 156820 97060 157020 97260
rect 156420 93060 156620 93260
rect 156020 93060 156220 93260
rect 155620 95860 155820 96060
rect 155620 92260 155820 92460
rect 156020 93460 156220 93660
rect 156420 97060 156620 97260
rect 155620 90660 155820 90860
rect 156020 90660 156220 90860
rect 156420 95060 156620 95260
rect 156820 95860 157020 96060
rect 156820 94660 157020 94860
rect 156420 95860 156620 96060
rect 155620 95060 155820 95260
rect 156820 94260 157020 94460
rect 156820 95060 157020 95260
rect 156420 92260 156620 92460
rect 155620 94660 155820 94860
rect 156820 95460 157020 95660
rect 155620 85860 155820 86060
rect 156020 89860 156220 90060
rect 156820 84660 157020 84860
rect 155620 85460 155820 85660
rect 156820 89860 157020 90060
rect 156020 89060 156220 89260
rect 156420 86660 156620 86860
rect 156420 85860 156620 86060
rect 156420 84660 156620 84860
rect 156820 86260 157020 86460
rect 156420 89460 156620 89660
rect 156820 89060 157020 89260
rect 155620 86260 155820 86460
rect 156420 86260 156620 86460
rect 155620 88260 155820 88460
rect 156820 85860 157020 86060
rect 156420 87060 156620 87260
rect 156420 85460 156620 85660
rect 156820 83860 157020 84060
rect 156420 83860 156620 84060
rect 155620 86660 155820 86860
rect 156420 87460 156620 87660
rect 155620 89860 155820 90060
rect 156020 83860 156220 84060
rect 156820 85460 157020 85660
rect 156020 87460 156220 87660
rect 156420 89860 156620 90060
rect 156420 87860 156620 88060
rect 155620 87060 155820 87260
rect 156820 86660 157020 86860
rect 156020 86260 156220 86460
rect 155620 88660 155820 88860
rect 156020 87860 156220 88060
rect 156020 88660 156220 88860
rect 155620 83860 155820 84060
rect 156820 87060 157020 87260
rect 156420 88260 156620 88460
rect 156020 85060 156220 85260
rect 156820 84260 157020 84460
rect 155620 87460 155820 87660
rect 156820 87460 157020 87660
rect 155620 84260 155820 84460
rect 156020 84260 156220 84460
rect 156420 84260 156620 84460
rect 156820 87860 157020 88060
rect 156020 85460 156220 85660
rect 156420 88660 156620 88860
rect 155620 84660 155820 84860
rect 156820 88260 157020 88460
rect 156820 85060 157020 85260
rect 156420 85060 156620 85260
rect 155620 87860 155820 88060
rect 155620 85060 155820 85260
rect 156820 88660 157020 88860
rect 155620 89460 155820 89660
rect 155620 89060 155820 89260
rect 156020 84660 156220 84860
rect 156020 85860 156220 86060
rect 156820 89460 157020 89660
rect 156020 89460 156220 89660
rect 156020 88260 156220 88460
rect 156020 86660 156220 86860
rect 156020 87060 156220 87260
rect 156420 89060 156620 89260
rect 156420 69460 156620 69660
rect 156020 69460 156220 69660
rect 156820 69460 157020 69660
rect 155620 69460 155820 69660
rect 156020 77860 156220 78060
rect 156820 79060 157020 79260
rect 156420 79060 156620 79260
rect 156820 79460 157020 79660
rect 156420 79460 156620 79660
rect 156820 79860 157020 80060
rect 156420 79860 156620 80060
rect 156020 78260 156220 78460
rect 156820 80260 157020 80460
rect 156420 80260 156620 80460
rect 156020 78660 156220 78860
rect 155620 77060 155820 77260
rect 156820 80660 157020 80860
rect 156420 80660 156620 80860
rect 156820 81060 157020 81260
rect 156420 81060 156620 81260
rect 156020 79060 156220 79260
rect 156820 81460 157020 81660
rect 156420 81460 156620 81660
rect 155620 79860 155820 80060
rect 156820 81860 157020 82060
rect 156420 81860 156620 82060
rect 156020 79460 156220 79660
rect 156820 82260 157020 82460
rect 156420 82260 156620 82460
rect 155620 78660 155820 78860
rect 155620 77460 155820 77660
rect 156020 79860 156220 80060
rect 156820 82660 157020 82860
rect 156420 82660 156620 82860
rect 156820 83060 157020 83260
rect 156420 83060 156620 83260
rect 155620 79460 155820 79660
rect 156020 80260 156220 80460
rect 156020 80660 156220 80860
rect 156020 81060 156220 81260
rect 155620 77860 155820 78060
rect 156820 78660 157020 78860
rect 156420 78660 156620 78860
rect 156020 83060 156220 83260
rect 155620 80660 155820 80860
rect 155620 81060 155820 81260
rect 156020 81860 156220 82060
rect 155620 81460 155820 81660
rect 155620 80260 155820 80460
rect 155620 79060 155820 79260
rect 156420 76660 156620 76860
rect 155620 81860 155820 82060
rect 156020 76660 156220 76860
rect 155620 82260 155820 82460
rect 156020 82260 156220 82460
rect 155620 82660 155820 82860
rect 156820 76660 157020 76860
rect 156420 77060 156620 77260
rect 156020 77060 156220 77260
rect 156820 77060 157020 77260
rect 155620 83060 155820 83260
rect 156820 77460 157020 77660
rect 155620 76660 155820 76860
rect 156820 77860 157020 78060
rect 156420 77860 156620 78060
rect 156020 82660 156220 82860
rect 156420 77460 156620 77660
rect 156020 77460 156220 77660
rect 156820 78260 157020 78460
rect 156420 78260 156620 78460
rect 156020 81460 156220 81660
rect 155620 78260 155820 78460
rect 156820 74260 157020 74460
rect 156020 74660 156220 74860
rect 156420 70260 156620 70460
rect 156420 76260 156620 76460
rect 156020 70260 156220 70460
rect 155620 74260 155820 74460
rect 156020 76260 156220 76460
rect 156420 73460 156620 73660
rect 156020 73460 156220 73660
rect 156420 71460 156620 71660
rect 156020 75860 156220 76060
rect 156420 70660 156620 70860
rect 156820 74660 157020 74860
rect 156020 70660 156220 70860
rect 156820 72660 157020 72860
rect 156020 71460 156220 71660
rect 155620 72260 155820 72460
rect 155620 71860 155820 72060
rect 155620 73060 155820 73260
rect 156420 71060 156620 71260
rect 156020 71060 156220 71260
rect 156820 75060 157020 75260
rect 155620 72660 155820 72860
rect 156820 73460 157020 73660
rect 155620 74660 155820 74860
rect 155620 71060 155820 71260
rect 155620 75460 155820 75660
rect 156020 75060 156220 75260
rect 156020 74260 156220 74460
rect 156020 75460 156220 75660
rect 156420 73860 156620 74060
rect 155620 70260 155820 70460
rect 156020 72260 156220 72460
rect 156820 75460 157020 75660
rect 156420 75860 156620 76060
rect 156420 72660 156620 72860
rect 156820 72260 157020 72460
rect 155620 75860 155820 76060
rect 155620 71460 155820 71660
rect 155620 69860 155820 70060
rect 156420 75460 156620 75660
rect 156020 72660 156220 72860
rect 156020 73860 156220 74060
rect 156820 71860 157020 72060
rect 156420 72260 156620 72460
rect 156820 70260 157020 70460
rect 156820 73860 157020 74060
rect 156820 73060 157020 73260
rect 156820 75860 157020 76060
rect 156420 73060 156620 73260
rect 155620 75060 155820 75260
rect 156420 71860 156620 72060
rect 156420 74260 156620 74460
rect 156420 69860 156620 70060
rect 156820 76260 157020 76460
rect 156820 71060 157020 71260
rect 155620 76260 155820 76460
rect 156020 71860 156220 72060
rect 156820 70660 157020 70860
rect 156020 69860 156220 70060
rect 156820 71460 157020 71660
rect 155620 73860 155820 74060
rect 156020 73060 156220 73260
rect 156820 69860 157020 70060
rect 156420 75060 156620 75260
rect 155620 70660 155820 70860
rect 155620 73460 155820 73660
rect 156420 74660 156620 74860
rect 156020 62660 156220 62860
rect 156820 62660 157020 62860
rect 156420 62660 156620 62860
rect 155620 62660 155820 62860
rect 156020 65460 156220 65660
rect 156020 68260 156220 68460
rect 156820 65860 157020 66060
rect 156820 66260 157020 66460
rect 155620 64660 155820 64860
rect 156020 65860 156220 66060
rect 156820 67060 157020 67260
rect 155620 66260 155820 66460
rect 156820 63860 157020 64060
rect 156420 64660 156620 64860
rect 156020 66260 156220 66460
rect 155620 68260 155820 68460
rect 156020 69060 156220 69260
rect 155620 69060 155820 69260
rect 156820 69060 157020 69260
rect 155620 65860 155820 66060
rect 156820 68260 157020 68460
rect 155620 65460 155820 65660
rect 156020 67060 156220 67260
rect 156020 63860 156220 64060
rect 156820 67860 157020 68060
rect 156420 68660 156620 68860
rect 156020 64260 156220 64460
rect 156420 67460 156620 67660
rect 156820 66660 157020 66860
rect 156820 64260 157020 64460
rect 156420 64260 156620 64460
rect 156820 68660 157020 68860
rect 156420 65060 156620 65260
rect 156420 67860 156620 68060
rect 156820 65060 157020 65260
rect 156420 63460 156620 63660
rect 156420 65460 156620 65660
rect 156020 68660 156220 68860
rect 155620 66660 155820 66860
rect 156020 67460 156220 67660
rect 156420 68260 156620 68460
rect 156420 63860 156620 64060
rect 156420 63060 156620 63260
rect 156420 65860 156620 66060
rect 155620 67460 155820 67660
rect 156020 66660 156220 66860
rect 156020 64660 156220 64860
rect 155620 64260 155820 64460
rect 155620 67060 155820 67260
rect 155620 63460 155820 63660
rect 156420 66260 156620 66460
rect 156820 65460 157020 65660
rect 156820 67460 157020 67660
rect 156820 64660 157020 64860
rect 156020 63460 156220 63660
rect 156020 65060 156220 65260
rect 155620 65060 155820 65260
rect 156420 66660 156620 66860
rect 155620 63860 155820 64060
rect 156020 63060 156220 63260
rect 156820 63060 157020 63260
rect 156420 67060 156620 67260
rect 155620 68660 155820 68860
rect 156020 67860 156220 68060
rect 155620 67860 155820 68060
rect 156820 63460 157020 63660
rect 155620 63060 155820 63260
rect 156420 69060 156620 69260
rect 156020 59060 156220 59260
rect 155620 59460 155820 59660
rect 156820 57460 157020 57660
rect 155620 56260 155820 56460
rect 155620 59860 155820 60060
rect 156420 57860 156620 58060
rect 156820 57860 157020 58060
rect 156420 60660 156620 60860
rect 155620 57460 155820 57660
rect 156020 61060 156220 61260
rect 156820 56260 157020 56460
rect 156420 56260 156620 56460
rect 156420 59460 156620 59660
rect 155620 60260 155820 60460
rect 156020 59460 156220 59660
rect 156820 60660 157020 60860
rect 156420 61460 156620 61660
rect 155620 56660 155820 56860
rect 156420 62260 156620 62460
rect 155620 61060 155820 61260
rect 156420 57060 156620 57260
rect 156820 61860 157020 62060
rect 156020 55860 156220 56060
rect 156820 59860 157020 60060
rect 156820 59460 157020 59660
rect 156020 56660 156220 56860
rect 156820 61460 157020 61660
rect 156820 56660 157020 56860
rect 156820 57060 157020 57260
rect 156420 61860 156620 62060
rect 156420 60260 156620 60460
rect 155620 61860 155820 62060
rect 155620 57860 155820 58060
rect 156420 59060 156620 59260
rect 156820 61060 157020 61260
rect 156020 58260 156220 58460
rect 156820 58660 157020 58860
rect 156420 59860 156620 60060
rect 156020 61460 156220 61660
rect 156420 55860 156620 56060
rect 156420 58260 156620 58460
rect 156020 62260 156220 62460
rect 155620 61460 155820 61660
rect 155620 55860 155820 56060
rect 155620 59060 155820 59260
rect 156020 59860 156220 60060
rect 156020 60660 156220 60860
rect 156420 61060 156620 61260
rect 156820 55860 157020 56060
rect 156420 56660 156620 56860
rect 156420 58660 156620 58860
rect 156020 58660 156220 58860
rect 156420 57460 156620 57660
rect 156820 59060 157020 59260
rect 156820 60260 157020 60460
rect 156020 57460 156220 57660
rect 156020 56260 156220 56460
rect 156820 62260 157020 62460
rect 156020 57060 156220 57260
rect 155620 60660 155820 60860
rect 156020 60260 156220 60460
rect 155620 57060 155820 57260
rect 156020 57860 156220 58060
rect 155620 58260 155820 58460
rect 156820 58260 157020 58460
rect 155620 62260 155820 62460
rect 156020 61860 156220 62060
rect 155620 58660 155820 58860
rect 700 83460 900 83660
rect 1100 83460 1300 83660
rect 1500 83460 1700 83660
rect 300 83460 500 83660
rect 1500 104260 1700 104460
rect 700 104260 900 104460
rect 1100 104260 1300 104460
rect 300 104260 500 104460
rect 1500 105860 1700 106060
rect 700 108260 900 108460
rect 1500 105460 1700 105660
rect 700 107860 900 108060
rect 1500 105060 1700 105260
rect 700 107460 900 107660
rect 1500 104660 1700 104860
rect 700 107060 900 107260
rect 1500 106660 1700 106860
rect 700 106660 900 106860
rect 700 106260 900 106460
rect 700 105860 900 106060
rect 700 105460 900 105660
rect 700 105060 900 105260
rect 700 104660 900 104860
rect 700 109060 900 109260
rect 1100 111060 1300 111260
rect 1100 110660 1300 110860
rect 1100 110260 1300 110460
rect 1100 109860 1300 110060
rect 1100 109460 1300 109660
rect 1100 109060 1300 109260
rect 1100 108660 1300 108860
rect 300 111060 500 111260
rect 1100 108260 1300 108460
rect 300 110660 500 110860
rect 1100 107860 1300 108060
rect 300 110260 500 110460
rect 1100 107460 1300 107660
rect 300 109860 500 110060
rect 1100 107060 1300 107260
rect 300 109460 500 109660
rect 1100 106660 1300 106860
rect 300 109060 500 109260
rect 1100 106260 1300 106460
rect 300 108660 500 108860
rect 700 109460 900 109660
rect 1100 105860 1300 106060
rect 300 108260 500 108460
rect 1100 105460 1300 105660
rect 300 107860 500 108060
rect 1100 105060 1300 105260
rect 300 107460 500 107660
rect 1100 104660 1300 104860
rect 300 107060 500 107260
rect 1500 106260 1700 106460
rect 300 106660 500 106860
rect 300 106260 500 106460
rect 300 105860 500 106060
rect 300 105460 500 105660
rect 300 105060 500 105260
rect 1500 111060 1700 111260
rect 300 104660 500 104860
rect 1500 110660 1700 110860
rect 700 108660 900 108860
rect 1500 110260 1700 110460
rect 1500 109860 1700 110060
rect 1500 109460 1700 109660
rect 1500 109060 1700 109260
rect 1500 108660 1700 108860
rect 700 111060 900 111260
rect 1500 108260 1700 108460
rect 700 110660 900 110860
rect 1500 107860 1700 108060
rect 700 110260 900 110460
rect 1500 107460 1700 107660
rect 700 109860 900 110060
rect 1500 107060 1700 107260
rect 700 98660 900 98860
rect 300 99060 500 99260
rect 1500 101860 1700 102060
rect 700 98260 900 98460
rect 1500 101460 1700 101660
rect 300 100260 500 100460
rect 700 97860 900 98060
rect 300 100660 500 100860
rect 1500 101060 1700 101260
rect 700 97460 900 97660
rect 700 103860 900 104060
rect 1500 100660 1700 100860
rect 700 103460 900 103660
rect 1500 100260 1700 100460
rect 700 103060 900 103260
rect 1500 99860 1700 100060
rect 1500 99460 1700 99660
rect 700 102660 900 102860
rect 1500 99060 1700 99260
rect 700 102260 900 102460
rect 300 97860 500 98060
rect 1500 98660 1700 98860
rect 700 101860 900 102060
rect 1100 103860 1300 104060
rect 300 99460 500 99660
rect 1100 103460 1300 103660
rect 1500 98260 1700 98460
rect 1100 103060 1300 103260
rect 700 101460 900 101660
rect 1100 102660 1300 102860
rect 1500 97860 1700 98060
rect 1100 102260 1300 102460
rect 1500 103860 1700 104060
rect 1500 97460 1700 97660
rect 1100 101860 1300 102060
rect 700 101060 900 101260
rect 300 97460 500 97660
rect 1100 101460 1300 101660
rect 700 100660 900 100860
rect 1100 97860 1300 98060
rect 300 103860 500 104060
rect 1100 101060 1300 101260
rect 300 98660 500 98860
rect 300 103460 500 103660
rect 1100 100660 1300 100860
rect 700 100260 900 100460
rect 300 103060 500 103260
rect 1100 100260 1300 100460
rect 1500 103460 1700 103660
rect 300 102660 500 102860
rect 1100 99860 1300 100060
rect 700 99860 900 100060
rect 300 102260 500 102460
rect 300 99860 500 100060
rect 1100 99460 1300 99660
rect 1500 103060 1700 103260
rect 300 101860 500 102060
rect 700 99460 900 99660
rect 1100 99060 1300 99260
rect 1100 97460 1300 97660
rect 300 101460 500 101660
rect 1500 102660 1700 102860
rect 1100 98660 1300 98860
rect 700 99060 900 99260
rect 300 101060 500 101260
rect 300 98260 500 98460
rect 1100 98260 1300 98460
rect 1500 102260 1700 102460
rect 1100 90260 1300 90460
rect 1500 90260 1700 90460
rect 700 90260 900 90460
rect 300 90260 500 90460
rect 1100 91460 1300 91660
rect 1500 93860 1700 94060
rect 300 97060 500 97260
rect 1500 93460 1700 93660
rect 300 94260 500 94460
rect 1100 91060 1300 91260
rect 1500 93060 1700 93260
rect 1100 90660 1300 90860
rect 300 93860 500 94060
rect 1500 92660 1700 92860
rect 1100 94260 1300 94460
rect 700 97060 900 97260
rect 1100 91860 1300 92060
rect 1500 92260 1700 92460
rect 300 96660 500 96860
rect 700 96660 900 96860
rect 1500 91860 1700 92060
rect 300 93460 500 93660
rect 1500 91460 1700 91660
rect 700 96260 900 96460
rect 1500 91060 1700 91260
rect 700 95860 900 96060
rect 1100 93860 1300 94060
rect 1500 90660 1700 90860
rect 300 93060 500 93260
rect 700 95460 900 95660
rect 1100 95460 1300 95660
rect 1100 94660 1300 94860
rect 700 95060 900 95260
rect 300 96260 500 96460
rect 700 94660 900 94860
rect 300 92660 500 92860
rect 700 94260 900 94460
rect 1100 96260 1300 96460
rect 1100 93460 1300 93660
rect 700 93860 900 94060
rect 1100 97060 1300 97260
rect 700 93460 900 93660
rect 300 92260 500 92460
rect 300 95860 500 96060
rect 700 93060 900 93260
rect 1100 93060 1300 93260
rect 1500 97060 1700 97260
rect 700 92660 900 92860
rect 300 91860 500 92060
rect 1100 96660 1300 96860
rect 700 92260 900 92460
rect 1500 96660 1700 96860
rect 300 91460 500 91660
rect 700 91860 900 92060
rect 1100 92660 1300 92860
rect 1500 96260 1700 96460
rect 700 91460 900 91660
rect 300 91060 500 91260
rect 300 95460 500 95660
rect 700 91060 900 91260
rect 1500 95860 1700 96060
rect 1100 95060 1300 95260
rect 700 90660 900 90860
rect 300 90660 500 90860
rect 1500 95460 1700 95660
rect 300 94660 500 94860
rect 1100 92260 1300 92460
rect 1500 95060 1700 95260
rect 1500 94260 1700 94460
rect 300 95060 500 95260
rect 1100 95860 1300 96060
rect 1500 94660 1700 94860
rect 300 89060 500 89260
rect 300 89460 500 89660
rect 1500 88660 1700 88860
rect 300 85060 500 85260
rect 300 87860 500 88060
rect 1100 85060 1300 85260
rect 1500 85060 1700 85260
rect 1500 88260 1700 88460
rect 300 84660 500 84860
rect 1100 88660 1300 88860
rect 700 85460 900 85660
rect 1500 87860 1700 88060
rect 1100 84260 1300 84460
rect 700 84260 900 84460
rect 300 84260 500 84460
rect 1500 87460 1700 87660
rect 300 87460 500 87660
rect 1500 84260 1700 84460
rect 700 85060 900 85260
rect 1100 88260 1300 88460
rect 1500 87060 1700 87260
rect 300 83860 500 84060
rect 700 88660 900 88860
rect 700 87860 900 88060
rect 300 88660 500 88860
rect 700 86260 900 86460
rect 1500 86660 1700 86860
rect 300 87060 500 87260
rect 1100 87860 1300 88060
rect 1100 89860 1300 90060
rect 700 87460 900 87660
rect 1500 85460 1700 85660
rect 700 83860 900 84060
rect 300 89860 500 90060
rect 1100 87460 1300 87660
rect 300 86660 500 86860
rect 1100 83860 1300 84060
rect 1500 83860 1700 84060
rect 1100 85460 1300 85660
rect 1100 87060 1300 87260
rect 300 88260 500 88460
rect 300 86260 500 86460
rect 1100 89460 1300 89660
rect 1100 84660 1300 84860
rect 1100 86660 1300 86860
rect 1500 89860 1700 90060
rect 1500 84660 1700 84860
rect 300 85860 500 86060
rect 700 87060 900 87260
rect 700 88260 900 88460
rect 1500 89460 1700 89660
rect 700 84660 900 84860
rect 1100 86260 1300 86460
rect 1500 86260 1700 86460
rect 700 89060 900 89260
rect 700 89860 900 90060
rect 700 86660 900 86860
rect 700 85860 900 86060
rect 1500 89060 1700 89260
rect 300 85460 500 85660
rect 700 89460 900 89660
rect 1100 85860 1300 86060
rect 1500 85860 1700 86060
rect 1100 89060 1300 89260
rect 300 69460 500 69660
rect 1500 69460 1700 69660
rect 700 69460 900 69660
rect 1100 69460 1300 69660
rect 300 77860 500 78060
rect 700 81060 900 81260
rect 700 80660 900 80860
rect 700 80260 900 80460
rect 300 79460 500 79660
rect 1100 83060 1300 83260
rect 1500 83060 1700 83260
rect 1100 82660 1300 82860
rect 1500 82660 1700 82860
rect 700 79860 900 80060
rect 300 77460 500 77660
rect 300 78660 500 78860
rect 1100 82260 1300 82460
rect 1500 82260 1700 82460
rect 700 79460 900 79660
rect 1100 81860 1300 82060
rect 1500 81860 1700 82060
rect 300 79860 500 80060
rect 1100 81460 1300 81660
rect 1500 81460 1700 81660
rect 700 79060 900 79260
rect 1100 81060 1300 81260
rect 1500 81060 1700 81260
rect 1100 80660 1300 80860
rect 1500 80660 1700 80860
rect 300 77060 500 77260
rect 700 78660 900 78860
rect 1100 80260 1300 80460
rect 1500 80260 1700 80460
rect 700 78260 900 78460
rect 1100 79860 1300 80060
rect 1500 79860 1700 80060
rect 1100 79460 1300 79660
rect 1500 79460 1700 79660
rect 1100 79060 1300 79260
rect 1500 79060 1700 79260
rect 700 77860 900 78060
rect 700 83060 900 83260
rect 1100 78660 1300 78860
rect 1500 78660 1700 78860
rect 300 78260 500 78460
rect 700 81460 900 81660
rect 1100 78260 1300 78460
rect 1500 78260 1700 78460
rect 700 77460 900 77660
rect 1100 77460 1300 77660
rect 700 82660 900 82860
rect 1100 77860 1300 78060
rect 1500 77860 1700 78060
rect 300 76660 500 76860
rect 1500 77460 1700 77660
rect 300 83060 500 83260
rect 1500 77060 1700 77260
rect 700 77060 900 77260
rect 1100 77060 1300 77260
rect 1500 76660 1700 76860
rect 300 82660 500 82860
rect 700 82260 900 82460
rect 300 82260 500 82460
rect 700 76660 900 76860
rect 300 81860 500 82060
rect 1100 76660 1300 76860
rect 300 79060 500 79260
rect 300 80260 500 80460
rect 300 81460 500 81660
rect 700 81860 900 82060
rect 300 81060 500 81260
rect 300 80660 500 80860
rect 300 71060 500 71260
rect 1500 73460 1700 73660
rect 300 72660 500 72860
rect 700 71060 900 71260
rect 1100 71060 1300 71260
rect 300 71860 500 72060
rect 300 72260 500 72460
rect 1500 72660 1700 72860
rect 700 70660 900 70860
rect 1100 70660 1300 70860
rect 700 75860 900 76060
rect 700 73460 900 73660
rect 1100 73460 1300 73660
rect 300 74260 500 74460
rect 700 70260 900 70460
rect 1100 70260 1300 70460
rect 700 74660 900 74860
rect 1100 74660 1300 74860
rect 300 70660 500 70860
rect 700 73060 900 73260
rect 700 69860 900 70060
rect 1100 69860 1300 70060
rect 1100 73060 1300 73260
rect 1500 71860 1700 72060
rect 300 71460 500 71660
rect 1100 75860 1300 76060
rect 700 75460 900 75660
rect 300 73860 500 74060
rect 300 75060 500 75260
rect 700 72660 900 72860
rect 1100 72660 1300 72860
rect 700 74260 900 74460
rect 1100 74260 1300 74460
rect 1100 75460 1300 75660
rect 300 70260 500 70460
rect 1500 73060 1700 73260
rect 700 72260 900 72460
rect 1100 72260 1300 72460
rect 1500 70660 1700 70860
rect 300 75860 500 76060
rect 300 75460 500 75660
rect 1500 71060 1700 71260
rect 300 73460 500 73660
rect 1500 69860 1700 70060
rect 1500 71460 1700 71660
rect 700 71860 900 72060
rect 1500 76260 1700 76460
rect 1100 71860 1300 72060
rect 1500 75860 1700 76060
rect 1500 70260 1700 70460
rect 700 73860 900 74060
rect 300 69860 500 70060
rect 1500 72260 1700 72460
rect 1500 75460 1700 75660
rect 1100 73860 1300 74060
rect 700 75060 900 75260
rect 300 74660 500 74860
rect 1500 75060 1700 75260
rect 300 73060 500 73260
rect 700 71460 900 71660
rect 1500 74660 1700 74860
rect 1100 71460 1300 71660
rect 700 76260 900 76460
rect 1100 76260 1300 76460
rect 1500 74260 1700 74460
rect 1100 75060 1300 75260
rect 300 76260 500 76460
rect 1500 73860 1700 74060
rect 1100 62660 1300 62860
rect 1500 62660 1700 62860
rect 300 62660 500 62860
rect 700 62660 900 62860
rect 300 65860 500 66060
rect 1500 66660 1700 66860
rect 1100 64660 1300 64860
rect 700 65860 900 66060
rect 1500 67460 1700 67660
rect 1500 63060 1700 63260
rect 300 64260 500 64460
rect 1100 63460 1300 63660
rect 700 64260 900 64460
rect 700 67060 900 67260
rect 300 69060 500 69260
rect 1500 63860 1700 64060
rect 1500 66260 1700 66460
rect 300 63860 500 64060
rect 300 68660 500 68860
rect 700 68660 900 68860
rect 700 63860 900 64060
rect 300 64660 500 64860
rect 1500 67860 1700 68060
rect 300 65460 500 65660
rect 700 65460 900 65660
rect 700 69060 900 69260
rect 1100 69060 1300 69260
rect 1100 63060 1300 63260
rect 1100 68660 1300 68860
rect 300 68260 500 68460
rect 700 68260 900 68460
rect 300 63460 500 63660
rect 1500 69060 1700 69260
rect 1500 65860 1700 66060
rect 1100 68260 1300 68460
rect 700 63460 900 63660
rect 1500 68260 1700 68460
rect 300 66260 500 66460
rect 1500 63460 1700 63660
rect 1100 67860 1300 68060
rect 1500 67060 1700 67260
rect 700 66260 900 66460
rect 1100 67460 1300 67660
rect 1500 64260 1700 64460
rect 300 63060 500 63260
rect 300 67860 500 68060
rect 700 67860 900 68060
rect 1100 67060 1300 67260
rect 700 63060 900 63260
rect 1100 66660 1300 66860
rect 300 65060 500 65260
rect 700 65060 900 65260
rect 1500 64660 1700 64860
rect 1500 65460 1700 65660
rect 1100 66260 1300 66460
rect 300 67060 500 67260
rect 700 64660 900 64860
rect 700 66660 900 66860
rect 300 67460 500 67660
rect 1100 65860 1300 66060
rect 1100 63860 1300 64060
rect 700 67460 900 67660
rect 300 66660 500 66860
rect 1100 65460 1300 65660
rect 1500 65060 1700 65260
rect 1100 65060 1300 65260
rect 1500 68660 1700 68860
rect 1100 64260 1300 64460
rect 1100 62260 1300 62460
rect 1100 61460 1300 61660
rect 700 59460 900 59660
rect 1100 59460 1300 59660
rect 1500 56260 1700 56460
rect 300 57460 500 57660
rect 1500 57860 1700 58060
rect 300 59860 500 60060
rect 1500 57460 1700 57660
rect 700 59060 900 59260
rect 700 61860 900 62060
rect 1500 58260 1700 58460
rect 300 57060 500 57260
rect 300 60660 500 60860
rect 1500 62260 1700 62460
rect 1500 60260 1700 60460
rect 700 58660 900 58860
rect 1100 56660 1300 56860
rect 700 60660 900 60860
rect 300 59060 500 59260
rect 300 61460 500 61660
rect 700 61460 900 61660
rect 700 58260 900 58460
rect 1100 59060 1300 59260
rect 1100 61860 1300 62060
rect 1500 61460 1700 61660
rect 700 55860 900 56060
rect 300 56660 500 56860
rect 300 56260 500 56460
rect 700 57860 900 58060
rect 1100 58660 1300 58860
rect 1100 58260 1300 58460
rect 1500 56660 1700 56860
rect 300 60260 500 60460
rect 700 60260 900 60460
rect 1100 60260 1300 60460
rect 300 57860 500 58060
rect 300 58260 500 58460
rect 700 57460 900 57660
rect 1100 61060 1300 61260
rect 1100 55860 1300 56060
rect 300 61860 500 62060
rect 1500 59860 1700 60060
rect 1500 60660 1700 60860
rect 1100 60660 1300 60860
rect 300 58660 500 58860
rect 700 57060 900 57260
rect 1500 55860 1700 56060
rect 1500 58660 1700 58860
rect 1500 57060 1700 57260
rect 1100 57060 1300 57260
rect 300 59460 500 59660
rect 700 59860 900 60060
rect 700 56660 900 56860
rect 300 55860 500 56060
rect 1100 56260 1300 56460
rect 1500 59060 1700 59260
rect 1100 59860 1300 60060
rect 1500 61860 1700 62060
rect 1100 57860 1300 58060
rect 700 56260 900 56460
rect 1500 61060 1700 61260
rect 1500 59460 1700 59660
rect 1100 57460 1300 57660
rect 300 61060 500 61260
rect 300 62260 500 62460
rect 700 62260 900 62460
rect 700 61060 900 61260
rect 300 27860 500 28060
rect 1100 27860 1300 28060
rect 1500 27860 1700 28060
rect 700 27860 900 28060
rect 700 41860 900 42060
rect 300 41860 500 42060
rect 1100 41860 1300 42060
rect 1500 41860 1700 42060
rect 700 48660 900 48860
rect 1100 48660 1300 48860
rect 300 48660 500 48860
rect 1500 48660 1700 48860
rect 1100 50260 1300 50460
rect 700 54660 900 54860
rect 1100 51060 1300 51260
rect 1100 49860 1300 50060
rect 700 52660 900 52860
rect 1100 49460 1300 49660
rect 1100 49060 1300 49260
rect 1100 50660 1300 50860
rect 700 52260 900 52460
rect 700 54260 900 54460
rect 300 55460 500 55660
rect 700 51860 900 52060
rect 300 55060 500 55260
rect 1100 55460 1300 55660
rect 300 54660 500 54860
rect 1100 55060 1300 55260
rect 1500 55460 1700 55660
rect 300 54260 500 54460
rect 1500 55060 1700 55260
rect 300 53860 500 54060
rect 700 51460 900 51660
rect 1100 54660 1300 54860
rect 1500 54660 1700 54860
rect 300 53460 500 53660
rect 1100 54260 1300 54460
rect 1500 54260 1700 54460
rect 300 53060 500 53260
rect 1500 53860 1700 54060
rect 300 52660 500 52860
rect 700 51060 900 51260
rect 1100 53860 1300 54060
rect 1500 53460 1700 53660
rect 700 53860 900 54060
rect 300 52260 500 52460
rect 1100 53460 1300 53660
rect 1500 53060 1700 53260
rect 300 51860 500 52060
rect 1500 52660 1700 52860
rect 300 51460 500 51660
rect 700 55060 900 55260
rect 1100 53060 1300 53260
rect 700 50660 900 50860
rect 1500 52260 1700 52460
rect 300 51060 500 51260
rect 1500 51860 1700 52060
rect 1100 52660 1300 52860
rect 300 50660 500 50860
rect 1500 51460 1700 51660
rect 300 50260 500 50460
rect 1500 51060 1700 51260
rect 300 49860 500 50060
rect 1100 52260 1300 52460
rect 1500 50660 1700 50860
rect 300 49460 500 49660
rect 700 50260 900 50460
rect 1500 50260 1700 50460
rect 300 49060 500 49260
rect 700 53460 900 53660
rect 700 49460 900 49660
rect 1500 49860 1700 50060
rect 1100 51860 1300 52060
rect 700 55460 900 55660
rect 1500 49460 1700 49660
rect 700 49860 900 50060
rect 1500 49060 1700 49260
rect 1100 51460 1300 51660
rect 700 49060 900 49260
rect 700 53060 900 53260
rect 1100 47060 1300 47260
rect 1500 47460 1700 47660
rect 1500 46660 1700 46860
rect 700 44660 900 44860
rect 1100 44260 1300 44460
rect 700 46260 900 46460
rect 1500 43860 1700 44060
rect 700 42260 900 42460
rect 1100 46660 1300 46860
rect 1500 43060 1700 43260
rect 1100 43860 1300 44060
rect 300 44260 500 44460
rect 700 44260 900 44460
rect 1500 45060 1700 45260
rect 1500 47860 1700 48060
rect 700 47460 900 47660
rect 300 46260 500 46460
rect 300 42660 500 42860
rect 1100 43460 1300 43660
rect 1100 48260 1300 48460
rect 1100 46260 1300 46460
rect 300 46660 500 46860
rect 700 43860 900 44060
rect 1100 43060 1300 43260
rect 700 45860 900 46060
rect 300 45460 500 45660
rect 1500 44260 1700 44460
rect 1500 45860 1700 46060
rect 1100 42660 1300 42860
rect 700 47060 900 47260
rect 1500 42660 1700 42860
rect 1100 47860 1300 48060
rect 1100 42260 1300 42460
rect 700 43460 900 43660
rect 1100 45860 1300 46060
rect 1500 46260 1700 46460
rect 300 43860 500 44060
rect 300 45860 500 46060
rect 300 43060 500 43260
rect 700 45460 900 45660
rect 1100 45460 1300 45660
rect 300 44660 500 44860
rect 1500 44660 1700 44860
rect 1100 47460 1300 47660
rect 700 43060 900 43260
rect 1500 43460 1700 43660
rect 700 47860 900 48060
rect 1500 42260 1700 42460
rect 300 45060 500 45260
rect 300 42260 500 42460
rect 1100 45060 1300 45260
rect 700 45060 900 45260
rect 300 48260 500 48460
rect 700 46660 900 46860
rect 300 43460 500 43660
rect 700 42660 900 42860
rect 300 47860 500 48060
rect 700 48260 900 48460
rect 300 47060 500 47260
rect 300 47460 500 47660
rect 1500 47060 1700 47260
rect 1100 44660 1300 44860
rect 1500 45460 1700 45660
rect 1500 48260 1700 48460
rect 700 36660 900 36860
rect 300 38660 500 38860
rect 700 39460 900 39660
rect 1500 37460 1700 37660
rect 700 36260 900 36460
rect 1100 35460 1300 35660
rect 300 36260 500 36460
rect 1500 39460 1700 39660
rect 300 38260 500 38460
rect 700 41060 900 41260
rect 700 35860 900 36060
rect 700 39060 900 39260
rect 1500 37060 1700 37260
rect 300 35860 500 36060
rect 700 35460 900 35660
rect 1500 40660 1700 40860
rect 1100 36260 1300 36460
rect 1500 39060 1700 39260
rect 700 38660 900 38860
rect 300 37860 500 38060
rect 1500 36660 1700 36860
rect 700 35060 900 35260
rect 300 35460 500 35660
rect 300 39460 500 39660
rect 700 40660 900 40860
rect 1100 37060 1300 37260
rect 700 38260 900 38460
rect 1500 36260 1700 36460
rect 300 35060 500 35260
rect 1100 39060 1300 39260
rect 1100 35060 1300 35260
rect 1500 38660 1700 38860
rect 1100 37860 1300 38060
rect 300 37460 500 37660
rect 1500 35860 1700 36060
rect 1100 35860 1300 36060
rect 700 37860 900 38060
rect 1100 37460 1300 37660
rect 300 41460 500 41660
rect 1100 38660 1300 38860
rect 1500 40260 1700 40460
rect 700 40260 900 40460
rect 1100 38260 1300 38460
rect 300 39060 500 39260
rect 1500 35460 1700 35660
rect 700 41460 900 41660
rect 1500 38260 1700 38460
rect 1100 41460 1300 41660
rect 1500 41060 1700 41260
rect 300 37060 500 37260
rect 1100 41060 1300 41260
rect 700 37460 900 37660
rect 300 40260 500 40460
rect 1500 41460 1700 41660
rect 1100 40660 1300 40860
rect 300 41060 500 41260
rect 700 39860 900 40060
rect 1500 35060 1700 35260
rect 1500 39860 1700 40060
rect 1100 40260 1300 40460
rect 700 37060 900 37260
rect 1500 37860 1700 38060
rect 1100 36660 1300 36860
rect 300 39860 500 40060
rect 1100 39860 1300 40060
rect 300 36660 500 36860
rect 1100 39460 1300 39660
rect 300 40660 500 40860
rect 1100 30660 1300 30860
rect 700 30260 900 30460
rect 700 33860 900 34060
rect 1100 31460 1300 31660
rect 300 29060 500 29260
rect 1500 34660 1700 34860
rect 1500 32260 1700 32460
rect 300 29860 500 30060
rect 1500 31860 1700 32060
rect 1500 29060 1700 29260
rect 300 34660 500 34860
rect 700 33460 900 33660
rect 1100 32660 1300 32860
rect 300 30260 500 30460
rect 300 31460 500 31660
rect 1500 31060 1700 31260
rect 300 33060 500 33260
rect 1100 29460 1300 29660
rect 700 33060 900 33260
rect 700 29060 900 29260
rect 300 32260 500 32460
rect 1500 33060 1700 33260
rect 1100 28260 1300 28460
rect 300 31860 500 32060
rect 1500 33460 1700 33660
rect 700 32660 900 32860
rect 300 30660 500 30860
rect 300 34260 500 34460
rect 1500 29460 1700 29660
rect 300 29460 500 29660
rect 1100 33460 1300 33660
rect 300 28660 500 28860
rect 700 32260 900 32460
rect 1500 28660 1700 28860
rect 300 32660 500 32860
rect 1100 29860 1300 30060
rect 700 34660 900 34860
rect 1100 31060 1300 31260
rect 300 31060 500 31260
rect 1500 30660 1700 30860
rect 1500 29860 1700 30060
rect 700 31860 900 32060
rect 1100 31860 1300 32060
rect 1500 31460 1700 31660
rect 300 28260 500 28460
rect 700 29860 900 30060
rect 300 33860 500 34060
rect 700 29460 900 29660
rect 700 31460 900 31660
rect 700 28660 900 28860
rect 1100 28660 1300 28860
rect 1100 29060 1300 29260
rect 1100 30260 1300 30460
rect 700 34260 900 34460
rect 1500 28260 1700 28460
rect 700 31060 900 31260
rect 1100 33060 1300 33260
rect 700 28260 900 28460
rect 1100 32260 1300 32460
rect 1500 32660 1700 32860
rect 1100 34660 1300 34860
rect 1500 33860 1700 34060
rect 1100 34260 1300 34460
rect 700 30660 900 30860
rect 1500 34260 1700 34460
rect 1100 33860 1300 34060
rect 300 33460 500 33660
rect 1500 30260 1700 30460
rect 1100 21060 1300 21260
rect 1500 21060 1700 21260
rect 700 21060 900 21260
rect 300 21060 500 21260
rect 1100 24660 1300 24860
rect 300 27460 500 27660
rect 1500 21460 1700 21660
rect 1500 23860 1700 24060
rect 300 27060 500 27260
rect 700 21460 900 21660
rect 700 25460 900 25660
rect 1100 23060 1300 23260
rect 300 26660 500 26860
rect 700 27060 900 27260
rect 700 22660 900 22860
rect 1500 23460 1700 23660
rect 300 26260 500 26460
rect 1500 25060 1700 25260
rect 300 21460 500 21660
rect 1100 23460 1300 23660
rect 700 26260 900 26460
rect 300 25860 500 26060
rect 1500 21860 1700 22060
rect 1100 27460 1300 27660
rect 1100 22660 1300 22860
rect 700 25060 900 25260
rect 1100 25460 1300 25660
rect 1100 25060 1300 25260
rect 1100 24260 1300 24460
rect 300 25460 500 25660
rect 1500 24660 1700 24860
rect 700 27460 900 27660
rect 300 25060 500 25260
rect 1100 27060 1300 27260
rect 700 23860 900 24060
rect 300 24660 500 24860
rect 1100 22260 1300 22460
rect 700 22260 900 22460
rect 1500 27460 1700 27660
rect 300 24260 500 24460
rect 1500 22660 1700 22860
rect 1100 26660 1300 26860
rect 300 23860 500 24060
rect 1500 27060 1700 27260
rect 700 23060 900 23260
rect 1100 23860 1300 24060
rect 700 24660 900 24860
rect 1500 22260 1700 22460
rect 300 23460 500 23660
rect 1500 26660 1700 26860
rect 1100 21860 1300 22060
rect 300 23060 500 23260
rect 1500 26260 1700 26460
rect 1100 26260 1300 26460
rect 700 23460 900 23660
rect 300 22660 500 22860
rect 700 26660 900 26860
rect 700 25860 900 26060
rect 700 24260 900 24460
rect 1500 25860 1700 26060
rect 300 22260 500 22460
rect 700 21860 900 22060
rect 1500 23060 1700 23260
rect 300 21860 500 22060
rect 1500 25460 1700 25660
rect 1100 21460 1300 21660
rect 1500 24260 1700 24460
rect 1100 25860 1300 26060
rect 300 14260 500 14460
rect 700 20660 900 20860
rect 300 16660 500 16860
rect 1100 14660 1300 14860
rect 700 19460 900 19660
rect 1100 18660 1300 18860
rect 1500 18660 1700 18860
rect 1100 15860 1300 16060
rect 700 17860 900 18060
rect 1500 15860 1700 16060
rect 300 15860 500 16060
rect 300 18660 500 18860
rect 700 19860 900 20060
rect 1500 15060 1700 15260
rect 1500 19860 1700 20060
rect 1500 20660 1700 20860
rect 700 15060 900 15260
rect 1100 18260 1300 18460
rect 300 14660 500 14860
rect 1100 19860 1300 20060
rect 700 18660 900 18860
rect 300 17860 500 18060
rect 1100 20660 1300 20860
rect 700 14260 900 14460
rect 300 16260 500 16460
rect 300 17060 500 17260
rect 300 19060 500 19260
rect 1500 16660 1700 16860
rect 700 15460 900 15660
rect 1100 17860 1300 18060
rect 1100 15460 1300 15660
rect 1500 19060 1700 19260
rect 1500 16260 1700 16460
rect 300 20660 500 20860
rect 700 17460 900 17660
rect 300 20260 500 20460
rect 300 19860 500 20060
rect 1100 17460 1300 17660
rect 1100 14260 1300 14460
rect 700 20260 900 20460
rect 1500 18260 1700 18460
rect 1500 17060 1700 17260
rect 300 19460 500 19660
rect 300 18260 500 18460
rect 1500 14660 1700 14860
rect 300 15460 500 15660
rect 700 16660 900 16860
rect 700 19060 900 19260
rect 1100 19460 1300 19660
rect 1500 19460 1700 19660
rect 1100 17060 1300 17260
rect 700 18260 900 18460
rect 1500 15460 1700 15660
rect 1100 16260 1300 16460
rect 1500 20260 1700 20460
rect 1100 20260 1300 20460
rect 300 17460 500 17660
rect 1100 16660 1300 16860
rect 1100 15060 1300 15260
rect 700 16260 900 16460
rect 1500 17460 1700 17660
rect 1100 19060 1300 19260
rect 700 17060 900 17260
rect 700 15860 900 16060
rect 700 14660 900 14860
rect 300 15060 500 15260
rect 1500 17860 1700 18060
rect 1500 14260 1700 14460
rect 1500 7060 1700 7260
rect 1100 7060 1300 7260
rect 300 7060 500 7260
rect 700 7060 900 7260
rect 1100 9860 1300 10060
rect 700 13460 900 13660
rect 1100 11860 1300 12060
rect 1500 8660 1700 8860
rect 300 7860 500 8060
rect 300 9060 500 9260
rect 300 7460 500 7660
rect 700 9860 900 10060
rect 1500 10660 1700 10860
rect 1100 7860 1300 8060
rect 300 10660 500 10860
rect 1100 13060 1300 13260
rect 1100 13460 1300 13660
rect 1100 11060 1300 11260
rect 1500 11860 1700 12060
rect 300 12260 500 12460
rect 1500 7460 1700 7660
rect 700 9460 900 9660
rect 700 11860 900 12060
rect 300 9860 500 10060
rect 700 11060 900 11260
rect 1500 9460 1700 9660
rect 1500 8260 1700 8460
rect 1500 12260 1700 12460
rect 700 9060 900 9260
rect 1500 13060 1700 13260
rect 700 13060 900 13260
rect 1500 9060 1700 9260
rect 700 13860 900 14060
rect 1100 7460 1300 7660
rect 300 11460 500 11660
rect 300 8660 500 8860
rect 1100 8260 1300 8460
rect 1500 10260 1700 10460
rect 300 13860 500 14060
rect 700 8660 900 8860
rect 300 13460 500 13660
rect 1500 11060 1700 11260
rect 1100 10260 1300 10460
rect 700 12260 900 12460
rect 700 10660 900 10860
rect 1100 10660 1300 10860
rect 300 9460 500 9660
rect 1100 11460 1300 11660
rect 300 13060 500 13260
rect 1500 12660 1700 12860
rect 700 8260 900 8460
rect 1100 9060 1300 9260
rect 1500 7860 1700 8060
rect 1100 12660 1300 12860
rect 1500 13460 1700 13660
rect 300 12660 500 12860
rect 700 12660 900 12860
rect 300 8260 500 8460
rect 700 7860 900 8060
rect 1500 13860 1700 14060
rect 1100 12260 1300 12460
rect 1100 9460 1300 9660
rect 1100 8660 1300 8860
rect 300 10260 500 10460
rect 1500 11460 1700 11660
rect 1500 9860 1700 10060
rect 300 11860 500 12060
rect 1100 13860 1300 14060
rect 700 10260 900 10460
rect 300 11060 500 11260
rect 700 7460 900 7660
rect 700 11460 900 11660
rect 1500 1460 1700 1660
rect 300 3060 500 3260
rect 700 2260 900 2460
rect 700 5860 900 6060
rect 1500 4260 1700 4460
rect 1100 3860 1300 4060
rect 300 2260 500 2460
rect 1100 5860 1300 6060
rect 700 2660 900 2860
rect 1500 660 1700 860
rect 700 3460 900 3660
rect 1500 5860 1700 6060
rect 1100 2660 1300 2860
rect 1100 3460 1300 3660
rect 300 1860 500 2060
rect 700 4660 900 4860
rect 700 6260 900 6460
rect 700 6660 900 6860
rect 1500 6660 1700 6860
rect 300 1060 500 1260
rect 300 5060 500 5260
rect 300 6660 500 6860
rect 1100 260 1300 460
rect 1500 2260 1700 2460
rect 700 660 900 860
rect 300 5460 500 5660
rect 300 6260 500 6460
rect 1500 2660 1700 2860
rect 300 4260 500 4460
rect 700 1460 900 1660
rect 1100 660 1300 860
rect 1500 5460 1700 5660
rect 700 260 900 460
rect 300 3860 500 4060
rect 1100 6660 1300 6860
rect 700 3860 900 4060
rect 1500 1060 1700 1260
rect 300 260 500 460
rect 700 1060 900 1260
rect 1500 3860 1700 4060
rect 1500 3060 1700 3260
rect 700 1860 900 2060
rect 700 5460 900 5660
rect 1100 1060 1300 1260
rect 700 3060 900 3260
rect 300 5860 500 6060
rect 1100 1860 1300 2060
rect 1100 5060 1300 5260
rect 1100 6260 1300 6460
rect 1100 4660 1300 4860
rect 700 4260 900 4460
rect 1500 5060 1700 5260
rect 300 2660 500 2860
rect 1500 6260 1700 6460
rect 1500 1860 1700 2060
rect 1500 4660 1700 4860
rect 1100 1460 1300 1660
rect 1500 3460 1700 3660
rect 300 1460 500 1660
rect 1100 5460 1300 5660
rect 1100 4260 1300 4460
rect 300 4660 500 4860
rect 300 660 500 860
rect 1100 3060 1300 3260
rect 1500 260 1700 460
rect 300 3460 500 3660
rect 700 5060 900 5260
rect 1100 2260 1300 2460
rect 156020 27860 156220 28060
rect 156820 27860 157020 28060
rect 156420 27860 156620 28060
rect 155620 27860 155820 28060
rect 156820 41860 157020 42060
rect 156420 41860 156620 42060
rect 155620 41860 155820 42060
rect 156020 41860 156220 42060
rect 156820 48660 157020 48860
rect 155620 48660 155820 48860
rect 156420 48660 156620 48860
rect 156020 48660 156220 48860
rect 156020 52260 156220 52460
rect 156420 50660 156620 50860
rect 156420 49060 156620 49260
rect 156420 49460 156620 49660
rect 156020 52660 156220 52860
rect 156420 49860 156620 50060
rect 156420 51060 156620 51260
rect 156020 54660 156220 54860
rect 156420 50260 156620 50460
rect 155620 55060 155820 55260
rect 156020 51860 156220 52060
rect 155620 55460 155820 55660
rect 156020 54260 156220 54460
rect 155620 54660 155820 54860
rect 156420 55460 156620 55660
rect 156820 55460 157020 55660
rect 156420 55060 156620 55260
rect 156020 53060 156220 53260
rect 156020 49060 156220 49260
rect 156420 51460 156620 51660
rect 156820 49060 157020 49260
rect 156020 49860 156220 50060
rect 156820 49460 157020 49660
rect 156020 55460 156220 55660
rect 156420 51860 156620 52060
rect 156820 49860 157020 50060
rect 156020 49460 156220 49660
rect 156020 53460 156220 53660
rect 155620 49060 155820 49260
rect 156820 50260 157020 50460
rect 156020 50260 156220 50460
rect 155620 49460 155820 49660
rect 156820 50660 157020 50860
rect 156420 52260 156620 52460
rect 155620 49860 155820 50060
rect 156820 51060 157020 51260
rect 155620 50260 155820 50460
rect 156820 51460 157020 51660
rect 155620 50660 155820 50860
rect 156420 52660 156620 52860
rect 156820 51860 157020 52060
rect 155620 51060 155820 51260
rect 156820 52260 157020 52460
rect 156020 50660 156220 50860
rect 156420 53060 156620 53260
rect 156020 55060 156220 55260
rect 155620 51460 155820 51660
rect 156820 52660 157020 52860
rect 155620 51860 155820 52060
rect 156820 53060 157020 53260
rect 156420 53460 156620 53660
rect 155620 52260 155820 52460
rect 156020 53860 156220 54060
rect 156820 53460 157020 53660
rect 156420 53860 156620 54060
rect 156020 51060 156220 51260
rect 155620 52660 155820 52860
rect 156820 53860 157020 54060
rect 155620 53060 155820 53260
rect 156820 54260 157020 54460
rect 156420 54260 156620 54460
rect 155620 53460 155820 53660
rect 156820 54660 157020 54860
rect 156420 54660 156620 54860
rect 156020 51460 156220 51660
rect 155620 53860 155820 54060
rect 156820 55060 157020 55260
rect 155620 54260 155820 54460
rect 156420 45860 156620 46060
rect 156820 42260 157020 42460
rect 156020 44660 156220 44860
rect 156020 43460 156220 43660
rect 156420 47460 156620 47660
rect 155620 47060 155820 47260
rect 156420 46660 156620 46860
rect 156420 42260 156620 42460
rect 156820 46660 157020 46860
rect 156020 47460 156220 47660
rect 156420 47860 156620 48060
rect 156820 48260 157020 48460
rect 156020 48260 156220 48460
rect 156820 47460 157020 47660
rect 156820 42660 157020 42860
rect 156820 44660 157020 44860
rect 156420 47060 156620 47260
rect 156020 47060 156220 47260
rect 155620 45060 155820 45260
rect 155620 47860 155820 48060
rect 155620 44660 155820 44860
rect 156420 42660 156620 42860
rect 156420 43860 156620 44060
rect 156820 45460 157020 45660
rect 156820 45860 157020 46060
rect 156020 42260 156220 42460
rect 156020 42660 156220 42860
rect 156420 45460 156620 45660
rect 156820 44260 157020 44460
rect 156820 45060 157020 45260
rect 156820 43460 157020 43660
rect 155620 45460 155820 45660
rect 156020 45460 156220 45660
rect 155620 43460 155820 43660
rect 155620 44260 155820 44460
rect 156020 45860 156220 46060
rect 156420 44660 156620 44860
rect 156820 43860 157020 44060
rect 156420 43060 156620 43260
rect 155620 43060 155820 43260
rect 156020 46660 156220 46860
rect 156820 43060 157020 43260
rect 156020 43860 156220 44060
rect 156020 44260 156220 44460
rect 155620 45860 155820 46060
rect 155620 46660 155820 46860
rect 156020 46260 156220 46460
rect 155620 48260 155820 48460
rect 156820 47060 157020 47260
rect 156420 46260 156620 46460
rect 155620 42260 155820 42460
rect 155620 43860 155820 44060
rect 156420 48260 156620 48460
rect 156020 43060 156220 43260
rect 156020 45060 156220 45260
rect 156020 47860 156220 48060
rect 156420 43460 156620 43660
rect 156820 46260 157020 46460
rect 156420 44260 156620 44460
rect 155620 42660 155820 42860
rect 155620 47460 155820 47660
rect 156420 45060 156620 45260
rect 156820 47860 157020 48060
rect 155620 46260 155820 46460
rect 155620 38660 155820 38860
rect 156020 41060 156220 41260
rect 155620 35860 155820 36060
rect 156020 36660 156220 36860
rect 155620 36260 155820 36460
rect 156020 35460 156220 35660
rect 156420 36260 156620 36460
rect 156020 39460 156220 39660
rect 155620 40660 155820 40860
rect 156420 39460 156620 39660
rect 156420 35460 156620 35660
rect 155620 36660 155820 36860
rect 156420 39860 156620 40060
rect 155620 39860 155820 40060
rect 156420 36660 156620 36860
rect 156820 37860 157020 38060
rect 156020 37060 156220 37260
rect 155620 38260 155820 38460
rect 156420 40260 156620 40460
rect 156820 39860 157020 40060
rect 156820 37060 157020 37260
rect 156820 35060 157020 35260
rect 156020 39860 156220 40060
rect 155620 41060 155820 41260
rect 156820 39060 157020 39260
rect 156420 40660 156620 40860
rect 156820 41460 157020 41660
rect 155620 40260 155820 40460
rect 156020 37460 156220 37660
rect 156420 41060 156620 41260
rect 155620 37060 155820 37260
rect 156020 35860 156220 36060
rect 156820 41060 157020 41260
rect 156020 36260 156220 36460
rect 156420 41460 156620 41660
rect 156820 38260 157020 38460
rect 156020 41460 156220 41660
rect 156820 35460 157020 35660
rect 156020 39060 156220 39260
rect 155620 39060 155820 39260
rect 156420 38260 156620 38460
rect 156020 40260 156220 40460
rect 156020 38660 156220 38860
rect 156820 40260 157020 40460
rect 156420 38660 156620 38860
rect 155620 41460 155820 41660
rect 155620 37860 155820 38060
rect 156420 37460 156620 37660
rect 156020 37860 156220 38060
rect 156420 35860 156620 36060
rect 156820 35860 157020 36060
rect 156820 40660 157020 40860
rect 155620 37460 155820 37660
rect 156420 37860 156620 38060
rect 156820 38660 157020 38860
rect 156420 35060 156620 35260
rect 156420 39060 156620 39260
rect 155620 35060 155820 35260
rect 156820 37460 157020 37660
rect 156820 36260 157020 36460
rect 156020 38260 156220 38460
rect 156420 37060 156620 37260
rect 156020 40660 156220 40860
rect 155620 39460 155820 39660
rect 156820 39460 157020 39660
rect 155620 35460 155820 35660
rect 156020 35060 156220 35260
rect 156820 36660 157020 36860
rect 155620 31060 155820 31260
rect 156420 29460 156620 29660
rect 155620 29460 155820 29660
rect 156820 29060 157020 29260
rect 156020 34260 156220 34460
rect 156820 31860 157020 32060
rect 156820 29460 157020 29660
rect 156420 29060 156620 29260
rect 156020 29460 156220 29660
rect 156420 31060 156620 31260
rect 155620 29860 155820 30060
rect 156820 30260 157020 30460
rect 156420 32260 156620 32460
rect 155620 34260 155820 34460
rect 156820 32260 157020 32460
rect 156020 34660 156220 34860
rect 156420 34260 156620 34460
rect 156820 34660 157020 34860
rect 155620 33060 155820 33260
rect 155620 29060 155820 29260
rect 155620 30660 155820 30860
rect 156420 29860 156620 30060
rect 155620 33860 155820 34060
rect 156820 32660 157020 32860
rect 156420 31460 156620 31660
rect 156420 28660 156620 28860
rect 156020 32660 156220 32860
rect 156020 33860 156220 34060
rect 155620 32660 155820 32860
rect 156020 31860 156220 32060
rect 156020 30260 156220 30460
rect 156820 33460 157020 33660
rect 156020 28260 156220 28460
rect 156020 31060 156220 31260
rect 156420 30660 156620 30860
rect 156820 28660 157020 28860
rect 156020 28660 156220 28860
rect 156820 31060 157020 31260
rect 156020 29860 156220 30060
rect 156020 32260 156220 32460
rect 155620 31860 155820 32060
rect 156020 33060 156220 33260
rect 155620 31460 155820 31660
rect 156420 31860 156620 32060
rect 156420 28260 156620 28460
rect 156820 34260 157020 34460
rect 156820 29860 157020 30060
rect 156420 34660 156620 34860
rect 156820 33860 157020 34060
rect 155620 28260 155820 28460
rect 155620 30260 155820 30460
rect 156820 33060 157020 33260
rect 155620 28660 155820 28860
rect 156420 33860 156620 34060
rect 156020 31460 156220 31660
rect 156420 32660 156620 32860
rect 156820 28260 157020 28460
rect 156420 33460 156620 33660
rect 155620 32260 155820 32460
rect 156420 30260 156620 30460
rect 156020 30660 156220 30860
rect 156820 30660 157020 30860
rect 156020 33460 156220 33660
rect 156420 33060 156620 33260
rect 155620 33460 155820 33660
rect 156020 29060 156220 29260
rect 155620 34660 155820 34860
rect 156820 31460 157020 31660
rect 156020 21060 156220 21260
rect 155620 21060 155820 21260
rect 156820 21060 157020 21260
rect 156420 21060 156620 21260
rect 155620 24660 155820 24860
rect 155620 22660 155820 22860
rect 156020 23860 156220 24060
rect 156420 27060 156620 27260
rect 156020 26660 156220 26860
rect 155620 25060 155820 25260
rect 156020 23460 156220 23660
rect 156020 27460 156220 27660
rect 156420 26260 156620 26460
rect 156820 24660 157020 24860
rect 156820 23060 157020 23260
rect 155620 25460 155820 25660
rect 156820 26260 157020 26460
rect 156420 24260 156620 24460
rect 156420 25060 156620 25260
rect 156420 25460 156620 25660
rect 155620 23060 155820 23260
rect 156820 24260 157020 24460
rect 156020 25060 156220 25260
rect 156420 22260 156620 22460
rect 156420 21860 156620 22060
rect 156420 22660 156620 22860
rect 156020 21860 156220 22060
rect 156420 27460 156620 27660
rect 156820 26660 157020 26860
rect 156820 21860 157020 22060
rect 155620 25860 155820 26060
rect 155620 23460 155820 23660
rect 156420 25860 156620 26060
rect 156020 26260 156220 26460
rect 156820 22260 157020 22460
rect 156420 23460 156620 23660
rect 155620 22260 155820 22460
rect 155620 21460 155820 21660
rect 156020 24660 156220 24860
rect 156420 21460 156620 21660
rect 156820 25060 157020 25260
rect 156420 23860 156620 24060
rect 155620 26260 155820 26460
rect 156820 23460 157020 23660
rect 156020 23060 156220 23260
rect 156820 25860 157020 26060
rect 156020 22660 156220 22860
rect 156820 27060 157020 27260
rect 156020 27060 156220 27260
rect 155620 26660 155820 26860
rect 155620 23860 155820 24060
rect 156420 23060 156620 23260
rect 155620 21860 155820 22060
rect 156420 26660 156620 26860
rect 156820 25460 157020 25660
rect 156020 25460 156220 25660
rect 156020 24260 156220 24460
rect 156020 21460 156220 21660
rect 156820 22660 157020 22860
rect 155620 27060 155820 27260
rect 156420 24660 156620 24860
rect 155620 24260 155820 24460
rect 156820 23860 157020 24060
rect 156820 21460 157020 21660
rect 156820 27460 157020 27660
rect 156020 25860 156220 26060
rect 155620 27460 155820 27660
rect 156020 22260 156220 22460
rect 156420 17460 156620 17660
rect 156820 17860 157020 18060
rect 155620 18660 155820 18860
rect 155620 15060 155820 15260
rect 155620 17060 155820 17260
rect 156020 15860 156220 16060
rect 156820 20660 157020 20860
rect 156820 15460 157020 15660
rect 156820 17060 157020 17260
rect 156420 15060 156620 15260
rect 156420 17060 156620 17260
rect 156420 19460 156620 19660
rect 155620 16660 155820 16860
rect 155620 15860 155820 16060
rect 155620 15460 155820 15660
rect 155620 18260 155820 18460
rect 155620 16260 155820 16460
rect 155620 17460 155820 17660
rect 156820 16660 157020 16860
rect 155620 14260 155820 14460
rect 156420 18260 156620 18460
rect 156820 15860 157020 16060
rect 156420 14660 156620 14860
rect 156820 19860 157020 20060
rect 155620 20260 155820 20460
rect 156020 17460 156220 17660
rect 156820 18260 157020 18460
rect 156420 17860 156620 18060
rect 156420 19060 156620 19260
rect 156020 17860 156220 18060
rect 156020 14260 156220 14460
rect 156420 16660 156620 16860
rect 156820 19060 157020 19260
rect 156020 20660 156220 20860
rect 156020 19060 156220 19260
rect 156820 19460 157020 19660
rect 156420 15860 156620 16060
rect 156820 14660 157020 14860
rect 156420 19860 156620 20060
rect 156820 15060 157020 15260
rect 155620 14660 155820 14860
rect 155620 19860 155820 20060
rect 156020 20260 156220 20460
rect 156420 20660 156620 20860
rect 156820 14260 157020 14460
rect 155620 19060 155820 19260
rect 155620 19460 155820 19660
rect 156820 18660 157020 18860
rect 156020 16260 156220 16460
rect 156420 16260 156620 16460
rect 156020 15460 156220 15660
rect 156420 20260 156620 20460
rect 156020 18260 156220 18460
rect 156820 16260 157020 16460
rect 156020 15060 156220 15260
rect 155620 17860 155820 18060
rect 156420 18660 156620 18860
rect 156020 17060 156220 17260
rect 156020 19860 156220 20060
rect 155620 20660 155820 20860
rect 156820 17460 157020 17660
rect 156420 14260 156620 14460
rect 156820 20260 157020 20460
rect 156020 18660 156220 18860
rect 156020 16660 156220 16860
rect 156420 15460 156620 15660
rect 156020 19460 156220 19660
rect 156020 14660 156220 14860
rect 156420 7060 156620 7260
rect 155620 7060 155820 7260
rect 156020 7060 156220 7260
rect 156820 7060 157020 7260
rect 156820 13860 157020 14060
rect 155620 8660 155820 8860
rect 156820 7860 157020 8060
rect 155620 11460 155820 11660
rect 155620 13860 155820 14060
rect 156420 7460 156620 7660
rect 155620 10260 155820 10460
rect 156020 13860 156220 14060
rect 156420 9060 156620 9260
rect 156820 9060 157020 9260
rect 156820 9860 157020 10060
rect 156020 13060 156220 13260
rect 156020 8260 156220 8460
rect 156820 13060 157020 13260
rect 156020 7860 156220 8060
rect 156020 9060 156220 9260
rect 156820 12660 157020 12860
rect 156420 12660 156620 12860
rect 156820 12260 157020 12460
rect 156420 8660 156620 8860
rect 156820 8260 157020 8460
rect 155620 13060 155820 13260
rect 156820 9460 157020 9660
rect 156020 11060 156220 11260
rect 155620 8260 155820 8460
rect 155620 9860 155820 10060
rect 156420 11460 156620 11660
rect 156020 11860 156220 12060
rect 156820 10260 157020 10460
rect 156020 9460 156220 9660
rect 156420 13860 156620 14060
rect 156820 7460 157020 7660
rect 155620 9460 155820 9660
rect 155620 12260 155820 12460
rect 155620 11860 155820 12060
rect 156820 11860 157020 12060
rect 156020 12660 156220 12860
rect 156420 10660 156620 10860
rect 156420 11060 156620 11260
rect 156420 13460 156620 13660
rect 156020 10660 156220 10860
rect 156420 8260 156620 8460
rect 156420 13060 156620 13260
rect 156420 9460 156620 9660
rect 155620 12660 155820 12860
rect 155620 10660 155820 10860
rect 156420 7860 156620 8060
rect 156020 12260 156220 12460
rect 156820 11460 157020 11660
rect 156820 10660 157020 10860
rect 156020 11460 156220 11660
rect 156420 10260 156620 10460
rect 156020 9860 156220 10060
rect 155620 7460 155820 7660
rect 156820 11060 157020 11260
rect 155620 9060 155820 9260
rect 156020 7460 156220 7660
rect 155620 7860 155820 8060
rect 156820 13460 157020 13660
rect 156820 8660 157020 8860
rect 155620 13460 155820 13660
rect 155620 11060 155820 11260
rect 156420 11860 156620 12060
rect 156020 13460 156220 13660
rect 156020 8660 156220 8860
rect 156420 12260 156620 12460
rect 156420 9860 156620 10060
rect 156020 10260 156220 10460
rect 156420 3460 156620 3660
rect 156020 2260 156220 2460
rect 155620 5460 155820 5660
rect 156420 5860 156620 6060
rect 155620 3860 155820 4060
rect 156420 3860 156620 4060
rect 155620 6660 155820 6860
rect 155620 1460 155820 1660
rect 155620 660 155820 860
rect 156820 260 157020 460
rect 156020 6660 156220 6860
rect 155620 3060 155820 3260
rect 156020 5460 156220 5660
rect 156820 5860 157020 6060
rect 156020 6260 156220 6460
rect 156020 260 156220 460
rect 155620 3460 155820 3660
rect 156420 260 156620 460
rect 156820 3460 157020 3660
rect 156420 5060 156620 5260
rect 156020 1060 156220 1260
rect 156420 4660 156620 4860
rect 156820 1460 157020 1660
rect 156820 6660 157020 6860
rect 156820 4260 157020 4460
rect 156020 660 156220 860
rect 156820 1060 157020 1260
rect 156420 1460 156620 1660
rect 155620 4660 155820 4860
rect 156020 2660 156220 2860
rect 156820 5060 157020 5260
rect 156020 4260 156220 4460
rect 155620 6260 155820 6460
rect 156020 3060 156220 3260
rect 156020 3460 156220 3660
rect 155620 1060 155820 1260
rect 155620 2260 155820 2460
rect 156020 1460 156220 1660
rect 156820 4660 157020 4860
rect 156420 1860 156620 2060
rect 156020 3860 156220 4060
rect 156420 1060 156620 1260
rect 156820 3860 157020 4060
rect 155620 260 155820 460
rect 156420 4260 156620 4460
rect 156820 2660 157020 2860
rect 156820 2260 157020 2460
rect 156820 1860 157020 2060
rect 156020 5860 156220 6060
rect 155620 5060 155820 5260
rect 156420 2260 156620 2460
rect 156420 2660 156620 2860
rect 156420 3060 156620 3260
rect 155620 1860 155820 2060
rect 155620 5860 155820 6060
rect 156420 660 156620 860
rect 156820 5460 157020 5660
rect 156820 660 157020 860
rect 156820 6260 157020 6460
rect 156020 4660 156220 4860
rect 156420 6260 156620 6460
rect 156820 3060 157020 3260
rect 156420 6660 156620 6860
rect 156020 1860 156220 2060
rect 156420 5460 156620 5660
rect 156020 5060 156220 5260
rect 155620 4260 155820 4460
rect 155620 2660 155820 2860
<< l69d44 >>
rect 84280 89527 84480 89727
rect 84280 89127 84480 89327
rect 84285 27472 84485 27672
rect 84285 27072 84485 27272
rect 156020 83460 156220 83660
rect 156420 83460 156620 83660
rect 156820 83460 157020 83660
rect 155620 83460 155820 83660
rect 156820 104260 157020 104460
rect 156020 104260 156220 104460
rect 156420 104260 156620 104460
rect 155620 104260 155820 104460
rect 156820 105860 157020 106060
rect 156020 108260 156220 108460
rect 156820 105460 157020 105660
rect 156020 107860 156220 108060
rect 156820 105060 157020 105260
rect 156020 107460 156220 107660
rect 156820 104660 157020 104860
rect 156020 107060 156220 107260
rect 156820 106660 157020 106860
rect 156020 106660 156220 106860
rect 156020 106260 156220 106460
rect 156020 105860 156220 106060
rect 156020 105460 156220 105660
rect 156020 105060 156220 105260
rect 156020 104660 156220 104860
rect 156020 109060 156220 109260
rect 156420 111060 156620 111260
rect 156420 110660 156620 110860
rect 156420 110260 156620 110460
rect 156420 109860 156620 110060
rect 156420 109460 156620 109660
rect 156420 109060 156620 109260
rect 156420 108660 156620 108860
rect 155620 111060 155820 111260
rect 156420 108260 156620 108460
rect 155620 110660 155820 110860
rect 156420 107860 156620 108060
rect 155620 110260 155820 110460
rect 156420 107460 156620 107660
rect 155620 109860 155820 110060
rect 156420 107060 156620 107260
rect 155620 109460 155820 109660
rect 156420 106660 156620 106860
rect 155620 109060 155820 109260
rect 156420 106260 156620 106460
rect 155620 108660 155820 108860
rect 156020 109460 156220 109660
rect 156420 105860 156620 106060
rect 155620 108260 155820 108460
rect 156420 105460 156620 105660
rect 155620 107860 155820 108060
rect 156420 105060 156620 105260
rect 155620 107460 155820 107660
rect 156420 104660 156620 104860
rect 155620 107060 155820 107260
rect 156820 106260 157020 106460
rect 155620 106660 155820 106860
rect 155620 106260 155820 106460
rect 155620 105860 155820 106060
rect 155620 105460 155820 105660
rect 155620 105060 155820 105260
rect 156820 111060 157020 111260
rect 155620 104660 155820 104860
rect 156820 110660 157020 110860
rect 156020 108660 156220 108860
rect 156820 110260 157020 110460
rect 156820 109860 157020 110060
rect 156820 109460 157020 109660
rect 156820 109060 157020 109260
rect 156820 108660 157020 108860
rect 156020 111060 156220 111260
rect 156820 108260 157020 108460
rect 156020 110660 156220 110860
rect 156820 107860 157020 108060
rect 156020 110260 156220 110460
rect 156820 107460 157020 107660
rect 156020 109860 156220 110060
rect 156820 107060 157020 107260
rect 156020 98660 156220 98860
rect 155620 99060 155820 99260
rect 156820 101860 157020 102060
rect 156020 98260 156220 98460
rect 156820 101460 157020 101660
rect 155620 100260 155820 100460
rect 156020 97860 156220 98060
rect 155620 100660 155820 100860
rect 156820 101060 157020 101260
rect 156020 97460 156220 97660
rect 156020 103860 156220 104060
rect 156820 100660 157020 100860
rect 156020 103460 156220 103660
rect 156820 100260 157020 100460
rect 156020 103060 156220 103260
rect 156820 99860 157020 100060
rect 156820 99460 157020 99660
rect 156020 102660 156220 102860
rect 156820 99060 157020 99260
rect 156020 102260 156220 102460
rect 155620 97860 155820 98060
rect 156820 98660 157020 98860
rect 156020 101860 156220 102060
rect 156420 103860 156620 104060
rect 155620 99460 155820 99660
rect 156420 103460 156620 103660
rect 156820 98260 157020 98460
rect 156420 103060 156620 103260
rect 156020 101460 156220 101660
rect 156420 102660 156620 102860
rect 156820 97860 157020 98060
rect 156420 102260 156620 102460
rect 156820 103860 157020 104060
rect 156820 97460 157020 97660
rect 156420 101860 156620 102060
rect 156020 101060 156220 101260
rect 155620 97460 155820 97660
rect 156420 101460 156620 101660
rect 156020 100660 156220 100860
rect 156420 97860 156620 98060
rect 155620 103860 155820 104060
rect 156420 101060 156620 101260
rect 155620 98660 155820 98860
rect 155620 103460 155820 103660
rect 156420 100660 156620 100860
rect 156020 100260 156220 100460
rect 155620 103060 155820 103260
rect 156420 100260 156620 100460
rect 156820 103460 157020 103660
rect 155620 102660 155820 102860
rect 156420 99860 156620 100060
rect 156020 99860 156220 100060
rect 155620 102260 155820 102460
rect 155620 99860 155820 100060
rect 156420 99460 156620 99660
rect 156820 103060 157020 103260
rect 155620 101860 155820 102060
rect 156020 99460 156220 99660
rect 156420 99060 156620 99260
rect 156420 97460 156620 97660
rect 155620 101460 155820 101660
rect 156820 102660 157020 102860
rect 156420 98660 156620 98860
rect 156020 99060 156220 99260
rect 155620 101060 155820 101260
rect 155620 98260 155820 98460
rect 156420 98260 156620 98460
rect 156820 102260 157020 102460
rect 156420 90260 156620 90460
rect 156820 90260 157020 90460
rect 156020 90260 156220 90460
rect 155620 90260 155820 90460
rect 156820 94260 157020 94460
rect 155620 95060 155820 95260
rect 156420 95860 156620 96060
rect 156820 94660 157020 94860
rect 156820 95460 157020 95660
rect 155620 94660 155820 94860
rect 156420 92260 156620 92460
rect 156820 95060 157020 95260
rect 156420 91460 156620 91660
rect 156820 93860 157020 94060
rect 155620 97060 155820 97260
rect 156820 93460 157020 93660
rect 155620 94260 155820 94460
rect 156420 91060 156620 91260
rect 156820 93060 157020 93260
rect 156420 90660 156620 90860
rect 155620 93860 155820 94060
rect 156820 92660 157020 92860
rect 156420 94260 156620 94460
rect 156020 97060 156220 97260
rect 156420 91860 156620 92060
rect 156820 92260 157020 92460
rect 155620 96660 155820 96860
rect 156020 96660 156220 96860
rect 156820 91860 157020 92060
rect 155620 93460 155820 93660
rect 156820 91460 157020 91660
rect 156020 96260 156220 96460
rect 156820 91060 157020 91260
rect 156020 95860 156220 96060
rect 156420 93860 156620 94060
rect 156820 90660 157020 90860
rect 155620 93060 155820 93260
rect 156020 95460 156220 95660
rect 156420 95460 156620 95660
rect 156420 94660 156620 94860
rect 156020 95060 156220 95260
rect 155620 96260 155820 96460
rect 156020 94660 156220 94860
rect 155620 92660 155820 92860
rect 156020 94260 156220 94460
rect 156420 96260 156620 96460
rect 156420 93460 156620 93660
rect 156020 93860 156220 94060
rect 156420 97060 156620 97260
rect 156020 93460 156220 93660
rect 155620 92260 155820 92460
rect 155620 95860 155820 96060
rect 156020 93060 156220 93260
rect 156420 93060 156620 93260
rect 156820 97060 157020 97260
rect 156020 92660 156220 92860
rect 155620 91860 155820 92060
rect 156420 96660 156620 96860
rect 156020 92260 156220 92460
rect 156820 96660 157020 96860
rect 155620 91460 155820 91660
rect 156020 91860 156220 92060
rect 156420 92660 156620 92860
rect 156820 96260 157020 96460
rect 156020 91460 156220 91660
rect 155620 91060 155820 91260
rect 155620 95460 155820 95660
rect 156020 91060 156220 91260
rect 156820 95860 157020 96060
rect 156420 95060 156620 95260
rect 156020 90660 156220 90860
rect 155620 90660 155820 90860
rect 155620 84660 155820 84860
rect 156020 86660 156220 86860
rect 156420 88660 156620 88860
rect 156020 85860 156220 86060
rect 156020 85460 156220 85660
rect 156820 89060 157020 89260
rect 156820 87860 157020 88060
rect 155620 85460 155820 85660
rect 156420 84260 156620 84460
rect 156020 89460 156220 89660
rect 156020 84260 156220 84460
rect 156420 85860 156620 86060
rect 155620 84260 155820 84460
rect 156820 85860 157020 86060
rect 156820 87460 157020 87660
rect 156420 89060 156620 89260
rect 155620 87460 155820 87660
rect 156820 84260 157020 84460
rect 156020 85060 156220 85260
rect 156420 88260 156620 88460
rect 156820 87060 157020 87260
rect 155620 83860 155820 84060
rect 156020 88660 156220 88860
rect 156020 87860 156220 88060
rect 155620 88660 155820 88860
rect 156020 86260 156220 86460
rect 156820 86660 157020 86860
rect 155620 87060 155820 87260
rect 156420 87860 156620 88060
rect 156420 89860 156620 90060
rect 156020 87460 156220 87660
rect 156820 85460 157020 85660
rect 156020 83860 156220 84060
rect 155620 89860 155820 90060
rect 156420 87460 156620 87660
rect 155620 86660 155820 86860
rect 156420 83860 156620 84060
rect 156820 83860 157020 84060
rect 156420 85460 156620 85660
rect 156420 87060 156620 87260
rect 155620 87860 155820 88060
rect 155620 88260 155820 88460
rect 156420 86260 156620 86460
rect 155620 86260 155820 86460
rect 156420 85060 156620 85260
rect 156420 89460 156620 89660
rect 156820 86260 157020 86460
rect 156420 84660 156620 84860
rect 156820 85060 157020 85260
rect 156420 86660 156620 86860
rect 156020 89060 156220 89260
rect 156820 89860 157020 90060
rect 156820 88260 157020 88460
rect 156820 84660 157020 84860
rect 156020 89860 156220 90060
rect 155620 85860 155820 86060
rect 155620 89060 155820 89260
rect 156020 87060 156220 87260
rect 155620 89460 155820 89660
rect 156020 88260 156220 88460
rect 156820 88660 157020 88860
rect 156820 89460 157020 89660
rect 155620 85060 155820 85260
rect 156020 84660 156220 84860
rect 107271 102067 107471 102267
rect 107721 102067 107921 102267
rect 108171 102067 108371 102267
rect 108621 102067 108821 102267
rect 109071 102067 109271 102267
rect 91267 103622 91467 103822
rect 91667 103622 91867 103822
rect 92067 103622 92267 103822
rect 92467 103622 92667 103822
rect 92867 103622 93067 103822
rect 93267 103622 93467 103822
rect 93667 103622 93867 103822
rect 94067 103622 94267 103822
rect 94467 103622 94667 103822
rect 94867 103622 95067 103822
rect 95267 103622 95467 103822
rect 95667 103622 95867 103822
rect 96067 103622 96267 103822
rect 96467 103622 96667 103822
rect 96867 103622 97067 103822
rect 97267 103622 97467 103822
rect 97667 103622 97867 103822
rect 98067 103622 98267 103822
rect 98467 103622 98667 103822
rect 98867 103622 99067 103822
rect 99267 103622 99467 103822
rect 99667 103622 99867 103822
rect 100067 103622 100267 103822
rect 100467 103622 100667 103822
rect 100867 103622 101067 103822
rect 101267 103622 101467 103822
rect 101667 103622 101867 103822
rect 102067 103622 102267 103822
rect 89267 103622 89467 103822
rect 89667 103622 89867 103822
rect 90067 103622 90267 103822
rect 90467 103622 90667 103822
rect 90867 103622 91067 103822
rect 85667 103622 85867 103822
rect 86067 103622 86267 103822
rect 86467 103622 86667 103822
rect 86867 103622 87067 103822
rect 87267 103622 87467 103822
rect 87667 103622 87867 103822
rect 88067 103622 88267 103822
rect 88467 103622 88667 103822
rect 88867 103622 89067 103822
rect 99815 86359 100015 86559
rect 99415 86359 99615 86559
rect 99815 86759 100015 86959
rect 99415 86759 99615 86959
rect 99815 87159 100015 87359
rect 99415 87159 99615 87359
rect 99815 87559 100015 87759
rect 99415 87559 99615 87759
rect 99815 87959 100015 88159
rect 99415 87959 99615 88159
rect 99815 88359 100015 88559
rect 99415 88359 99615 88559
rect 99815 88759 100015 88959
rect 99415 88759 99615 88959
rect 92280 89127 92480 89327
rect 91880 89527 92080 89727
rect 91880 89127 92080 89327
rect 91480 89527 91680 89727
rect 91480 89127 91680 89327
rect 91080 89527 91280 89727
rect 91080 89127 91280 89327
rect 90680 89527 90880 89727
rect 90680 89127 90880 89327
rect 90280 89527 90480 89727
rect 90280 89127 90480 89327
rect 89880 89527 90080 89727
rect 89880 89127 90080 89327
rect 89480 89527 89680 89727
rect 89480 89127 89680 89327
rect 89080 89527 89280 89727
rect 89080 89127 89280 89327
rect 88680 89527 88880 89727
rect 88680 89127 88880 89327
rect 88280 89527 88480 89727
rect 88280 89127 88480 89327
rect 87880 89527 88080 89727
rect 87880 89127 88080 89327
rect 87480 89527 87680 89727
rect 87480 89127 87680 89327
rect 87080 89527 87280 89727
rect 87080 89127 87280 89327
rect 86680 89527 86880 89727
rect 86680 89127 86880 89327
rect 86280 89527 86480 89727
rect 86280 89127 86480 89327
rect 85880 89527 86080 89727
rect 85880 89127 86080 89327
rect 85480 89527 85680 89727
rect 85480 89127 85680 89327
rect 85080 89527 85280 89727
rect 85080 89127 85280 89327
rect 84680 89527 84880 89727
rect 84680 89127 84880 89327
rect 99815 83559 100015 83759
rect 99415 83559 99615 83759
rect 96280 89527 96480 89727
rect 96280 89127 96480 89327
rect 95880 89527 96080 89727
rect 95880 89127 96080 89327
rect 95480 89527 95680 89727
rect 95480 89127 95680 89327
rect 95080 89527 95280 89727
rect 95080 89127 95280 89327
rect 94680 89527 94880 89727
rect 94680 89127 94880 89327
rect 94280 89527 94480 89727
rect 94280 89127 94480 89327
rect 93880 89527 94080 89727
rect 93880 89127 94080 89327
rect 93480 89527 93680 89727
rect 93480 89127 93680 89327
rect 93080 89527 93280 89727
rect 93080 89127 93280 89327
rect 92680 89527 92880 89727
rect 92680 89127 92880 89327
rect 92280 89527 92480 89727
rect 99815 83959 100015 84159
rect 99415 83959 99615 84159
rect 99815 84359 100015 84559
rect 99415 84359 99615 84559
rect 99815 84759 100015 84959
rect 99415 84759 99615 84959
rect 99815 85159 100015 85359
rect 99415 85159 99615 85359
rect 99815 85559 100015 85759
rect 99415 85559 99615 85759
rect 99815 85959 100015 86159
rect 99415 85959 99615 86159
rect 99815 69559 100015 69759
rect 99415 69559 99615 69759
rect 99815 74359 100015 74559
rect 99415 74359 99615 74559
rect 99815 74759 100015 74959
rect 99415 74759 99615 74959
rect 99815 75159 100015 75359
rect 99415 75159 99615 75359
rect 99815 75559 100015 75759
rect 99415 75559 99615 75759
rect 99815 75959 100015 76159
rect 99415 75959 99615 76159
rect 99815 76359 100015 76559
rect 99415 76359 99615 76559
rect 99815 76759 100015 76959
rect 99415 76759 99615 76959
rect 99815 77159 100015 77359
rect 99415 77159 99615 77359
rect 99815 77559 100015 77759
rect 99415 77559 99615 77759
rect 99815 77959 100015 78159
rect 99415 77959 99615 78159
rect 99815 78359 100015 78559
rect 99415 78359 99615 78559
rect 99815 78759 100015 78959
rect 99415 78759 99615 78959
rect 99815 79159 100015 79359
rect 99415 79159 99615 79359
rect 99815 79559 100015 79759
rect 99415 79559 99615 79759
rect 99815 79959 100015 80159
rect 99415 79959 99615 80159
rect 99815 80359 100015 80559
rect 99415 80359 99615 80559
rect 99815 80759 100015 80959
rect 99415 80759 99615 80959
rect 99815 81159 100015 81359
rect 99415 81159 99615 81359
rect 99815 81559 100015 81759
rect 99415 81559 99615 81759
rect 99815 81959 100015 82159
rect 99415 81959 99615 82159
rect 99815 82359 100015 82559
rect 99415 82359 99615 82559
rect 99815 82759 100015 82959
rect 99415 82759 99615 82959
rect 99815 83159 100015 83359
rect 99415 83159 99615 83359
rect 99815 73959 100015 74159
rect 99415 73959 99615 74159
rect 99815 69959 100015 70159
rect 99415 69959 99615 70159
rect 99815 70359 100015 70559
rect 99415 70359 99615 70559
rect 99815 70759 100015 70959
rect 99415 70759 99615 70959
rect 99815 71159 100015 71359
rect 99415 71159 99615 71359
rect 99815 71559 100015 71759
rect 99415 71559 99615 71759
rect 99815 71959 100015 72159
rect 99415 71959 99615 72159
rect 99815 72359 100015 72559
rect 99415 72359 99615 72559
rect 99815 72759 100015 72959
rect 99415 72759 99615 72959
rect 99815 73159 100015 73359
rect 99415 73159 99615 73359
rect 99815 73559 100015 73759
rect 99415 73559 99615 73759
rect 99415 61959 99615 62159
rect 99815 62359 100015 62559
rect 99415 62359 99615 62559
rect 99815 62759 100015 62959
rect 99415 62759 99615 62959
rect 99815 63159 100015 63359
rect 99415 63159 99615 63359
rect 99815 63559 100015 63759
rect 99415 63559 99615 63759
rect 99815 63959 100015 64159
rect 99415 63959 99615 64159
rect 99815 64359 100015 64559
rect 99415 64359 99615 64559
rect 99815 64759 100015 64959
rect 99415 64759 99615 64959
rect 99815 65159 100015 65359
rect 99415 65159 99615 65359
rect 99815 65559 100015 65759
rect 99815 55959 100015 56159
rect 99415 55959 99615 56159
rect 99815 56359 100015 56559
rect 99415 56359 99615 56559
rect 99815 56759 100015 56959
rect 99415 56759 99615 56959
rect 99815 57159 100015 57359
rect 99415 57159 99615 57359
rect 99815 57559 100015 57759
rect 99415 57559 99615 57759
rect 99815 57959 100015 58159
rect 99415 57959 99615 58159
rect 99815 58359 100015 58559
rect 99415 58359 99615 58559
rect 99815 58759 100015 58959
rect 99415 58759 99615 58959
rect 99815 59159 100015 59359
rect 99415 59159 99615 59359
rect 99815 59559 100015 59759
rect 99415 59559 99615 59759
rect 99815 59959 100015 60159
rect 99415 59959 99615 60159
rect 99815 60359 100015 60559
rect 99415 60359 99615 60559
rect 99815 60759 100015 60959
rect 99415 60759 99615 60959
rect 99815 69159 100015 69359
rect 99415 69159 99615 69359
rect 99815 61159 100015 61359
rect 99415 61159 99615 61359
rect 99815 61559 100015 61759
rect 99415 61559 99615 61759
rect 99815 61959 100015 62159
rect 99815 66759 100015 66959
rect 99415 66759 99615 66959
rect 99815 67159 100015 67359
rect 99415 67159 99615 67359
rect 99815 67559 100015 67759
rect 99415 67559 99615 67759
rect 99815 67959 100015 68159
rect 99415 67959 99615 68159
rect 99815 68359 100015 68559
rect 99415 68359 99615 68559
rect 99815 68759 100015 68959
rect 99415 68759 99615 68959
rect 99815 65959 100015 66159
rect 99415 65959 99615 66159
rect 99815 66359 100015 66559
rect 99415 66359 99615 66559
rect 99415 65559 99615 65759
rect 155620 69460 155820 69660
rect 156820 69460 157020 69660
rect 156020 69460 156220 69660
rect 156420 69460 156620 69660
rect 156020 82660 156220 82860
rect 156420 77860 156620 78060
rect 156820 77860 157020 78060
rect 155620 76660 155820 76860
rect 156820 77460 157020 77660
rect 155620 83060 155820 83260
rect 156820 77060 157020 77260
rect 156020 77060 156220 77260
rect 156420 77060 156620 77260
rect 156820 76660 157020 76860
rect 155620 82660 155820 82860
rect 156020 82260 156220 82460
rect 155620 82260 155820 82460
rect 156020 76660 156220 76860
rect 155620 81860 155820 82060
rect 156420 76660 156620 76860
rect 155620 79060 155820 79260
rect 155620 80260 155820 80460
rect 155620 81460 155820 81660
rect 156020 81860 156220 82060
rect 155620 81060 155820 81260
rect 155620 80660 155820 80860
rect 156420 78260 156620 78460
rect 156820 78260 157020 78460
rect 156020 77460 156220 77660
rect 156420 77460 156620 77660
rect 155620 77860 155820 78060
rect 156020 81060 156220 81260
rect 156020 80660 156220 80860
rect 156020 80260 156220 80460
rect 155620 79460 155820 79660
rect 156420 83060 156620 83260
rect 156820 83060 157020 83260
rect 156420 82660 156620 82860
rect 156820 82660 157020 82860
rect 156020 79860 156220 80060
rect 155620 77460 155820 77660
rect 155620 78660 155820 78860
rect 156420 82260 156620 82460
rect 156820 82260 157020 82460
rect 156020 79460 156220 79660
rect 156420 81860 156620 82060
rect 156820 81860 157020 82060
rect 155620 79860 155820 80060
rect 156420 81460 156620 81660
rect 156820 81460 157020 81660
rect 156020 79060 156220 79260
rect 156420 81060 156620 81260
rect 156820 81060 157020 81260
rect 156420 80660 156620 80860
rect 156820 80660 157020 80860
rect 155620 77060 155820 77260
rect 156020 78660 156220 78860
rect 156420 80260 156620 80460
rect 156820 80260 157020 80460
rect 156020 78260 156220 78460
rect 156420 79860 156620 80060
rect 156820 79860 157020 80060
rect 156420 79460 156620 79660
rect 156820 79460 157020 79660
rect 156420 79060 156620 79260
rect 156820 79060 157020 79260
rect 156020 77860 156220 78060
rect 156020 83060 156220 83260
rect 156420 78660 156620 78860
rect 156820 78660 157020 78860
rect 155620 78260 155820 78460
rect 156020 81460 156220 81660
rect 155620 70260 155820 70460
rect 156820 73060 157020 73260
rect 156020 72260 156220 72460
rect 156420 70660 156620 70860
rect 156420 72260 156620 72460
rect 156820 70660 157020 70860
rect 155620 75860 155820 76060
rect 155620 72660 155820 72860
rect 155620 75460 155820 75660
rect 156820 71060 157020 71260
rect 155620 73460 155820 73660
rect 156020 75860 156220 76060
rect 156820 69860 157020 70060
rect 156820 71460 157020 71660
rect 156020 71860 156220 72060
rect 156020 73460 156220 73660
rect 156820 76260 157020 76460
rect 156420 71860 156620 72060
rect 156820 75860 157020 76060
rect 156420 73460 156620 73660
rect 156820 70260 157020 70460
rect 156020 73860 156220 74060
rect 155620 69860 155820 70060
rect 156020 71060 156220 71260
rect 156820 72260 157020 72460
rect 156820 75460 157020 75660
rect 156420 73860 156620 74060
rect 155620 74260 155820 74460
rect 156020 75060 156220 75260
rect 155620 74660 155820 74860
rect 156820 75060 157020 75260
rect 156020 70260 156220 70460
rect 155620 73060 155820 73260
rect 156020 71460 156220 71660
rect 156820 74660 157020 74860
rect 156420 70260 156620 70460
rect 156420 71460 156620 71660
rect 156020 76260 156220 76460
rect 155620 71060 155820 71260
rect 156420 76260 156620 76460
rect 156820 74260 157020 74460
rect 156020 74660 156220 74860
rect 156420 75060 156620 75260
rect 155620 76260 155820 76460
rect 156420 74660 156620 74860
rect 156820 73860 157020 74060
rect 155620 70660 155820 70860
rect 156420 71060 156620 71260
rect 156020 73060 156220 73260
rect 156020 69860 156220 70060
rect 156420 69860 156620 70060
rect 155620 71860 155820 72060
rect 156420 73060 156620 73260
rect 156820 71860 157020 72060
rect 155620 71460 155820 71660
rect 155620 72260 155820 72460
rect 156420 75860 156620 76060
rect 156020 75460 156220 75660
rect 155620 73860 155820 74060
rect 156820 73460 157020 73660
rect 155620 75060 155820 75260
rect 156020 72660 156220 72860
rect 156420 72660 156620 72860
rect 156820 72660 157020 72860
rect 156020 74260 156220 74460
rect 156420 74260 156620 74460
rect 156420 75460 156620 75660
rect 156020 70660 156220 70860
rect 156420 62660 156620 62860
rect 156820 62660 157020 62860
rect 155620 62660 155820 62860
rect 156020 62660 156220 62860
rect 156020 65060 156220 65260
rect 156020 66660 156220 66860
rect 156420 66260 156620 66460
rect 156420 65860 156620 66060
rect 156820 68660 157020 68860
rect 155620 63060 155820 63260
rect 155620 67460 155820 67660
rect 155620 65060 155820 65260
rect 155620 67860 155820 68060
rect 156020 64660 156220 64860
rect 156420 66660 156620 66860
rect 155620 65860 155820 66060
rect 156820 66660 157020 66860
rect 156420 63860 156620 64060
rect 156420 64660 156620 64860
rect 156020 67860 156220 68060
rect 156020 65860 156220 66060
rect 156820 67460 157020 67660
rect 156820 63060 157020 63260
rect 155620 64260 155820 64460
rect 155620 67060 155820 67260
rect 156420 63460 156620 63660
rect 156820 64660 157020 64860
rect 156020 64260 156220 64460
rect 156420 67060 156620 67260
rect 156020 67060 156220 67260
rect 155620 69060 155820 69260
rect 156820 63860 157020 64060
rect 156820 66260 157020 66460
rect 155620 63860 155820 64060
rect 156020 67460 156220 67660
rect 155620 68660 155820 68860
rect 156020 68660 156220 68860
rect 156020 63860 156220 64060
rect 155620 64660 155820 64860
rect 156820 67860 157020 68060
rect 155620 65460 155820 65660
rect 156020 63060 156220 63260
rect 156020 65460 156220 65660
rect 156020 69060 156220 69260
rect 156420 69060 156620 69260
rect 156820 65060 157020 65260
rect 156420 63060 156620 63260
rect 156420 68660 156620 68860
rect 155620 68260 155820 68460
rect 155620 66660 155820 66860
rect 156020 68260 156220 68460
rect 155620 63460 155820 63660
rect 156820 69060 157020 69260
rect 156820 65860 157020 66060
rect 156420 68260 156620 68460
rect 156420 65060 156620 65260
rect 156020 63460 156220 63660
rect 156820 65460 157020 65660
rect 156820 68260 157020 68460
rect 155620 66260 155820 66460
rect 156820 63460 157020 63660
rect 156420 67860 156620 68060
rect 156820 67060 157020 67260
rect 156420 64260 156620 64460
rect 156020 66260 156220 66460
rect 156420 65460 156620 65660
rect 156420 67460 156620 67660
rect 156820 64260 157020 64460
rect 155620 60260 155820 60460
rect 156020 55860 156220 56060
rect 156020 62260 156220 62460
rect 156420 62260 156620 62460
rect 156820 57860 157020 58060
rect 155620 61460 155820 61660
rect 156820 60260 157020 60460
rect 156820 59060 157020 59260
rect 156020 61860 156220 62060
rect 156020 61060 156220 61260
rect 155620 59460 155820 59660
rect 156420 60660 156620 60860
rect 156020 60260 156220 60460
rect 156420 58660 156620 58860
rect 156820 59860 157020 60060
rect 156420 59060 156620 59260
rect 156820 57060 157020 57260
rect 156420 57460 156620 57660
rect 156420 61460 156620 61660
rect 156820 55860 157020 56060
rect 156820 58260 157020 58460
rect 156420 61860 156620 62060
rect 156020 56260 156220 56460
rect 156420 59860 156620 60060
rect 156420 60260 156620 60460
rect 155620 57460 155820 57660
rect 156020 58260 156220 58460
rect 155620 59860 155820 60060
rect 156420 59460 156620 59660
rect 156420 55860 156620 56060
rect 156820 56260 157020 56460
rect 156020 61460 156220 61660
rect 155620 57060 155820 57260
rect 156420 58260 156620 58460
rect 156420 57060 156620 57260
rect 156820 61860 157020 62060
rect 155620 57860 155820 58060
rect 156020 60660 156220 60860
rect 156020 57060 156220 57260
rect 156420 56660 156620 56860
rect 156820 59460 157020 59660
rect 155620 56660 155820 56860
rect 156020 59860 156220 60060
rect 155620 55860 155820 56060
rect 155620 60660 155820 60860
rect 156820 57460 157020 57660
rect 156820 61060 157020 61260
rect 155620 61060 155820 61260
rect 155620 58260 155820 58460
rect 156820 60660 157020 60860
rect 156020 57860 156220 58060
rect 156820 56660 157020 56860
rect 156020 59460 156220 59660
rect 155620 58660 155820 58860
rect 155620 56260 155820 56460
rect 156020 58660 156220 58860
rect 156820 62260 157020 62460
rect 156020 56660 156220 56860
rect 156820 61460 157020 61660
rect 155620 62260 155820 62460
rect 156020 57460 156220 57660
rect 156820 58660 157020 58860
rect 155620 59060 155820 59260
rect 156020 59060 156220 59260
rect 156420 56260 156620 56460
rect 156420 57860 156620 58060
rect 156420 61060 156620 61260
rect 155620 61860 155820 62060
rect 17138 83429 17338 83629
rect 16738 83429 16938 83629
rect 66280 89527 66480 89727
rect 66280 89127 66480 89327
rect 65880 89527 66080 89727
rect 65880 89127 66080 89327
rect 65480 89527 65680 89727
rect 65480 89127 65680 89327
rect 65080 89527 65280 89727
rect 65080 89127 65280 89327
rect 64680 89527 64880 89727
rect 64680 89127 64880 89327
rect 64280 89527 64480 89727
rect 64280 89127 64480 89327
rect 63880 89527 64080 89727
rect 63880 89127 64080 89327
rect 63480 89527 63680 89727
rect 63480 89127 63680 89327
rect 63080 89527 63280 89727
rect 63080 89127 63280 89327
rect 62680 89527 62880 89727
rect 62680 89127 62880 89327
rect 62280 89527 62480 89727
rect 62280 89127 62480 89327
rect 61880 89527 62080 89727
rect 61880 89127 62080 89327
rect 61480 89527 61680 89727
rect 61480 89127 61680 89327
rect 61080 89527 61280 89727
rect 61080 89127 61280 89327
rect 60680 89527 60880 89727
rect 60680 89127 60880 89327
rect 60280 89527 60480 89727
rect 60280 89127 60480 89327
rect 59880 89527 60080 89727
rect 59880 89127 60080 89327
rect 59480 89527 59680 89727
rect 59480 89127 59680 89327
rect 59080 89527 59280 89727
rect 59080 89127 59280 89327
rect 58680 89527 58880 89727
rect 58680 89127 58880 89327
rect 58280 89527 58480 89727
rect 58280 89127 58480 89327
rect 57880 89527 58080 89727
rect 57880 89127 58080 89327
rect 57480 89527 57680 89727
rect 57480 89127 57680 89327
rect 57080 89527 57280 89727
rect 57080 89127 57280 89327
rect 48270 91027 48470 91227
rect 48270 91427 48470 91627
rect 48670 91027 48870 91227
rect 48670 91427 48870 91627
rect 49070 91027 49270 91227
rect 49070 91427 49270 91627
rect 49470 91027 49670 91227
rect 49470 91427 49670 91627
rect 49870 91027 50070 91227
rect 49870 91427 50070 91627
rect 50270 91027 50470 91227
rect 50270 91427 50470 91627
rect 50670 91027 50870 91227
rect 50670 91427 50870 91627
rect 51070 91027 51270 91227
rect 51070 91427 51270 91627
rect 73480 89527 73680 89727
rect 73480 89127 73680 89327
rect 73080 89527 73280 89727
rect 73080 89127 73280 89327
rect 72680 89527 72880 89727
rect 72680 89127 72880 89327
rect 72280 89527 72480 89727
rect 72280 89127 72480 89327
rect 71880 89527 72080 89727
rect 71880 89127 72080 89327
rect 71480 89527 71680 89727
rect 71480 89127 71680 89327
rect 71080 89527 71280 89727
rect 71080 89127 71280 89327
rect 70680 89527 70880 89727
rect 70680 89127 70880 89327
rect 70280 89527 70480 89727
rect 70280 89127 70480 89327
rect 69880 89527 70080 89727
rect 69880 89127 70080 89327
rect 69480 89527 69680 89727
rect 69480 89127 69680 89327
rect 69080 89527 69280 89727
rect 69080 89127 69280 89327
rect 68680 89527 68880 89727
rect 68680 89127 68880 89327
rect 68280 89527 68480 89727
rect 68280 89127 68480 89327
rect 67880 89527 68080 89727
rect 67880 89127 68080 89327
rect 67480 89527 67680 89727
rect 67480 89127 67680 89327
rect 67080 89527 67280 89727
rect 67080 89127 67280 89327
rect 83880 89127 84080 89327
rect 83480 89527 83680 89727
rect 83480 89127 83680 89327
rect 83080 89527 83280 89727
rect 83080 89127 83280 89327
rect 82680 89527 82880 89727
rect 82680 89127 82880 89327
rect 82280 89527 82480 89727
rect 82280 89127 82480 89327
rect 81880 89527 82080 89727
rect 81880 89127 82080 89327
rect 81480 89527 81680 89727
rect 81480 89127 81680 89327
rect 81080 89527 81280 89727
rect 81080 89127 81280 89327
rect 80680 89527 80880 89727
rect 80680 89127 80880 89327
rect 80280 89527 80480 89727
rect 66680 89527 66880 89727
rect 66680 89127 66880 89327
rect 76280 89527 76480 89727
rect 76280 89127 76480 89327
rect 75880 89527 76080 89727
rect 75880 89127 76080 89327
rect 75480 89527 75680 89727
rect 75480 89127 75680 89327
rect 75080 89527 75280 89727
rect 75080 89127 75280 89327
rect 74680 89527 74880 89727
rect 74680 89127 74880 89327
rect 74280 89527 74480 89727
rect 74280 89127 74480 89327
rect 73880 89527 74080 89727
rect 73880 89127 74080 89327
rect 83880 89527 84080 89727
rect 79080 89527 79280 89727
rect 79080 89127 79280 89327
rect 78680 89527 78880 89727
rect 78680 89127 78880 89327
rect 78280 89527 78480 89727
rect 78280 89127 78480 89327
rect 77880 89527 78080 89727
rect 77880 89127 78080 89327
rect 77480 89527 77680 89727
rect 77480 89127 77680 89327
rect 77080 89527 77280 89727
rect 77080 89127 77280 89327
rect 79880 89527 80080 89727
rect 79880 89127 80080 89327
rect 79480 89527 79680 89727
rect 79480 89127 79680 89327
rect 80280 89127 80480 89327
rect 76680 89527 76880 89727
rect 76680 89127 76880 89327
rect 29870 91027 30070 91227
rect 29870 91427 30070 91627
rect 21070 91027 21270 91227
rect 21070 91427 21270 91627
rect 21470 91027 21670 91227
rect 21470 91427 21670 91627
rect 21870 91027 22070 91227
rect 21870 91427 22070 91627
rect 22270 91027 22470 91227
rect 22270 91427 22470 91627
rect 22670 91027 22870 91227
rect 22670 91427 22870 91627
rect 23070 91027 23270 91227
rect 23070 91427 23270 91627
rect 23470 91027 23670 91227
rect 23470 91427 23670 91627
rect 23870 91027 24070 91227
rect 23870 91427 24070 91627
rect 24270 91027 24470 91227
rect 24270 91427 24470 91627
rect 24670 91027 24870 91227
rect 24670 91427 24870 91627
rect 25070 91027 25270 91227
rect 25070 91427 25270 91627
rect 25470 91027 25670 91227
rect 25470 91427 25670 91627
rect 25870 91027 26070 91227
rect 25870 91427 26070 91627
rect 26270 91027 26470 91227
rect 26270 91427 26470 91627
rect 26670 91027 26870 91227
rect 26670 91427 26870 91627
rect 27070 91027 27270 91227
rect 27070 91427 27270 91627
rect 27470 91027 27670 91227
rect 27470 91427 27670 91627
rect 27870 91027 28070 91227
rect 28270 91027 28470 91227
rect 28270 91427 28470 91627
rect 28670 91027 28870 91227
rect 28670 91427 28870 91627
rect 29070 91027 29270 91227
rect 29070 91427 29270 91627
rect 29470 91027 29670 91227
rect 29470 91427 29670 91627
rect 27870 91427 28070 91627
rect 20670 91027 20870 91227
rect 20670 91427 20870 91627
rect 11870 91027 12070 91227
rect 11870 91427 12070 91627
rect 12270 91027 12470 91227
rect 12270 91427 12470 91627
rect 12670 91027 12870 91227
rect 12670 91427 12870 91627
rect 13070 91027 13270 91227
rect 13070 91427 13270 91627
rect 13470 91027 13670 91227
rect 13470 91427 13670 91627
rect 13870 91027 14070 91227
rect 13870 91427 14070 91627
rect 14270 91027 14470 91227
rect 14270 91427 14470 91627
rect 14670 91027 14870 91227
rect 14670 91427 14870 91627
rect 15070 91027 15270 91227
rect 15070 91427 15270 91627
rect 15470 91027 15670 91227
rect 15470 91427 15670 91627
rect 15870 91027 16070 91227
rect 15870 91427 16070 91627
rect 16270 91027 16470 91227
rect 16270 91427 16470 91627
rect 16670 91027 16870 91227
rect 16670 91427 16870 91627
rect 17070 91027 17270 91227
rect 17070 91427 17270 91627
rect 17470 91027 17670 91227
rect 17470 91427 17670 91627
rect 17870 91027 18070 91227
rect 17870 91427 18070 91627
rect 18270 91027 18470 91227
rect 18270 91427 18470 91627
rect 18670 91027 18870 91227
rect 18670 91427 18870 91627
rect 19070 91027 19270 91227
rect 19070 91427 19270 91627
rect 19470 91027 19670 91227
rect 19470 91427 19670 91627
rect 19870 91027 20070 91227
rect 19870 91427 20070 91627
rect 20270 91027 20470 91227
rect 20270 91427 20470 91627
rect 17138 87429 17338 87629
rect 16738 87429 16938 87629
rect 17138 87029 17338 87229
rect 17138 86629 17338 86829
rect 16738 86629 16938 86829
rect 16738 87029 16938 87229
rect 17138 83829 17338 84029
rect 16738 83829 16938 84029
rect 17138 84229 17338 84429
rect 16738 84229 16938 84429
rect 17138 84629 17338 84829
rect 16738 84629 16938 84829
rect 17138 85029 17338 85229
rect 16738 85029 16938 85229
rect 17138 85429 17338 85629
rect 16738 85429 16938 85629
rect 17138 85829 17338 86029
rect 16738 85829 16938 86029
rect 17138 86229 17338 86429
rect 16738 86229 16938 86429
rect 42270 91427 42470 91627
rect 42670 91027 42870 91227
rect 42670 91427 42870 91627
rect 30270 91027 30470 91227
rect 30270 91427 30470 91627
rect 30670 91027 30870 91227
rect 45070 91427 45270 91627
rect 30670 91427 30870 91627
rect 31070 91027 31270 91227
rect 31070 91427 31270 91627
rect 31470 91027 31670 91227
rect 31470 91427 31670 91627
rect 31870 91027 32070 91227
rect 31870 91427 32070 91627
rect 32270 91027 32470 91227
rect 32270 91427 32470 91627
rect 32670 91027 32870 91227
rect 32670 91427 32870 91627
rect 33070 91027 33270 91227
rect 33070 91427 33270 91627
rect 33470 91027 33670 91227
rect 33470 91427 33670 91627
rect 33870 91027 34070 91227
rect 33870 91427 34070 91627
rect 34270 91027 34470 91227
rect 45470 91027 45670 91227
rect 45470 91427 45670 91627
rect 45870 91027 46070 91227
rect 45870 91427 46070 91627
rect 46270 91027 46470 91227
rect 46270 91427 46470 91627
rect 46670 91027 46870 91227
rect 46670 91427 46870 91627
rect 47070 91027 47270 91227
rect 47070 91427 47270 91627
rect 47470 91027 47670 91227
rect 47470 91427 47670 91627
rect 47870 91027 48070 91227
rect 47870 91427 48070 91627
rect 34270 91427 34470 91627
rect 34670 91027 34870 91227
rect 34670 91427 34870 91627
rect 35070 91027 35270 91227
rect 35070 91427 35270 91627
rect 35470 91027 35670 91227
rect 35470 91427 35670 91627
rect 35870 91027 36070 91227
rect 35870 91427 36070 91627
rect 36270 91027 36470 91227
rect 36270 91427 36470 91627
rect 36670 91027 36870 91227
rect 36670 91427 36870 91627
rect 37070 91027 37270 91227
rect 37070 91427 37270 91627
rect 37470 91027 37670 91227
rect 43070 91027 43270 91227
rect 37470 91427 37670 91627
rect 37870 91027 38070 91227
rect 37870 91427 38070 91627
rect 38270 91027 38470 91227
rect 38270 91427 38470 91627
rect 38670 91027 38870 91227
rect 38670 91427 38870 91627
rect 39070 91027 39270 91227
rect 39070 91427 39270 91627
rect 39470 91027 39670 91227
rect 39470 91427 39670 91627
rect 39870 91027 40070 91227
rect 39870 91427 40070 91627
rect 40270 91027 40470 91227
rect 40270 91427 40470 91627
rect 40670 91027 40870 91227
rect 40670 91427 40870 91627
rect 41070 91027 41270 91227
rect 41070 91427 41270 91627
rect 41470 91027 41670 91227
rect 43070 91427 43270 91627
rect 43470 91027 43670 91227
rect 43470 91427 43670 91627
rect 43870 91027 44070 91227
rect 43870 91427 44070 91627
rect 44270 91027 44470 91227
rect 44270 91427 44470 91627
rect 44670 91027 44870 91227
rect 44670 91427 44870 91627
rect 45070 91027 45270 91227
rect 41470 91427 41670 91627
rect 41870 91027 42070 91227
rect 41870 91427 42070 91627
rect 42270 91027 42470 91227
rect 17138 69829 17338 70029
rect 16738 69829 16938 70029
rect 17138 70229 17338 70429
rect 16738 70229 16938 70429
rect 17138 70629 17338 70829
rect 16738 70629 16938 70829
rect 17138 71029 17338 71229
rect 16738 71029 16938 71229
rect 17138 71429 17338 71629
rect 16738 71429 16938 71629
rect 17138 71829 17338 72029
rect 16738 71829 16938 72029
rect 17138 72229 17338 72429
rect 16738 72229 16938 72429
rect 17138 72629 17338 72829
rect 16738 72629 16938 72829
rect 17138 73029 17338 73229
rect 16738 73029 16938 73229
rect 17138 73429 17338 73629
rect 16738 73429 16938 73629
rect 17138 73829 17338 74029
rect 16738 73829 16938 74029
rect 17138 74229 17338 74429
rect 16738 74229 16938 74429
rect 17138 74629 17338 74829
rect 16738 74629 16938 74829
rect 17138 75029 17338 75229
rect 16738 75029 16938 75229
rect 17138 75429 17338 75629
rect 16738 75429 16938 75629
rect 17138 75829 17338 76029
rect 16738 75829 16938 76029
rect 17138 76229 17338 76429
rect 16738 76229 16938 76429
rect 17138 76629 17338 76829
rect 16738 76629 16938 76829
rect 17138 77029 17338 77229
rect 16738 77029 16938 77229
rect 17138 77429 17338 77629
rect 16738 77429 16938 77629
rect 17138 77829 17338 78029
rect 16738 77829 16938 78029
rect 17138 78229 17338 78429
rect 16738 78229 16938 78429
rect 17138 78629 17338 78829
rect 16738 78629 16938 78829
rect 17138 79029 17338 79229
rect 16738 79029 16938 79229
rect 17138 79429 17338 79629
rect 16738 79429 16938 79629
rect 17138 79829 17338 80029
rect 16738 79829 16938 80029
rect 17138 80229 17338 80429
rect 16738 80229 16938 80429
rect 17138 80629 17338 80829
rect 16738 80629 16938 80829
rect 17138 81029 17338 81229
rect 16738 81029 16938 81229
rect 17138 81429 17338 81629
rect 16738 81429 16938 81629
rect 17138 81829 17338 82029
rect 16738 81829 16938 82029
rect 17138 82229 17338 82429
rect 16738 82229 16938 82429
rect 17138 82629 17338 82829
rect 16738 82629 16938 82829
rect 17138 83029 17338 83229
rect 16738 83029 16938 83229
rect 17138 66229 17338 66429
rect 16738 66229 16938 66429
rect 17138 66629 17338 66829
rect 16738 66629 16938 66829
rect 17138 67029 17338 67229
rect 16738 67029 16938 67229
rect 17138 67429 17338 67629
rect 16738 67429 16938 67629
rect 17138 64629 17338 64829
rect 16738 64629 16938 64829
rect 17138 65029 17338 65229
rect 16738 65029 16938 65229
rect 17138 67829 17338 68029
rect 16738 67829 16938 68029
rect 17138 68229 17338 68429
rect 16738 68229 16938 68429
rect 17138 68629 17338 68829
rect 16738 68629 16938 68829
rect 17138 69029 17338 69229
rect 16738 69029 16938 69229
rect 17138 69429 17338 69629
rect 16738 64229 16938 64429
rect 17138 55829 17338 56029
rect 16738 55829 16938 56029
rect 17138 56229 17338 56429
rect 16738 56229 16938 56429
rect 17138 56629 17338 56829
rect 16738 56629 16938 56829
rect 17138 57029 17338 57229
rect 16738 57029 16938 57229
rect 17138 57429 17338 57629
rect 16738 57429 16938 57629
rect 17138 57829 17338 58029
rect 16738 57829 16938 58029
rect 17138 58229 17338 58429
rect 16738 58229 16938 58429
rect 17138 58629 17338 58829
rect 16738 58629 16938 58829
rect 17138 59029 17338 59229
rect 16738 69429 16938 69629
rect 16738 62229 16938 62429
rect 17138 62629 17338 62829
rect 16738 62629 16938 62829
rect 17138 63029 17338 63229
rect 16738 63029 16938 63229
rect 17138 63429 17338 63629
rect 16738 63429 16938 63629
rect 17138 63829 17338 64029
rect 16738 63829 16938 64029
rect 17138 64229 17338 64429
rect 17138 65429 17338 65629
rect 16738 65429 16938 65629
rect 17138 65829 17338 66029
rect 16738 65829 16938 66029
rect 16738 59029 16938 59229
rect 17138 59429 17338 59629
rect 16738 59429 16938 59629
rect 17138 59829 17338 60029
rect 16738 59829 16938 60029
rect 17138 60229 17338 60429
rect 16738 60229 16938 60429
rect 17138 60629 17338 60829
rect 16738 60629 16938 60829
rect 17138 61029 17338 61229
rect 16738 61029 16938 61229
rect 17138 61429 17338 61629
rect 16738 61429 16938 61629
rect 17138 61829 17338 62029
rect 16738 61829 16938 62029
rect 17138 62229 17338 62429
rect 23188 27929 23388 28129
rect 22788 27929 22988 28129
rect 48090 17879 48290 18079
rect 48090 17479 48290 17679
rect 16738 49829 16938 50029
rect 17138 50229 17338 50429
rect 16738 50229 16938 50429
rect 17138 50629 17338 50829
rect 16738 50629 16938 50829
rect 17138 51029 17338 51229
rect 16738 51029 16938 51229
rect 17138 51429 17338 51629
rect 16738 51429 16938 51629
rect 17138 51829 17338 52029
rect 16738 51829 16938 52029
rect 17138 52229 17338 52429
rect 16738 52229 16938 52429
rect 17138 52629 17338 52829
rect 16738 52629 16938 52829
rect 17138 53029 17338 53229
rect 16738 53029 16938 53229
rect 17138 53429 17338 53629
rect 16738 53429 16938 53629
rect 17138 53829 17338 54029
rect 16738 53829 16938 54029
rect 17138 54229 17338 54429
rect 16738 54229 16938 54429
rect 17138 54629 17338 54829
rect 16738 54629 16938 54829
rect 17138 55029 17338 55229
rect 16738 55029 16938 55229
rect 17138 55429 17338 55629
rect 16738 55429 16938 55629
rect 17138 48229 17338 48429
rect 16738 48229 16938 48429
rect 17138 48629 17338 48829
rect 16738 48629 16938 48829
rect 17138 49029 17338 49229
rect 16738 49029 16938 49229
rect 17138 49429 17338 49629
rect 23188 41929 23388 42129
rect 22788 41929 22988 42129
rect 23188 42329 23388 42529
rect 22788 42329 22988 42529
rect 23188 42729 23388 42929
rect 22788 42729 22988 42929
rect 23188 43129 23388 43329
rect 22788 43129 22988 43329
rect 23188 43529 23388 43729
rect 22788 43529 22988 43729
rect 23188 43929 23388 44129
rect 22788 43929 22988 44129
rect 23188 44329 23388 44529
rect 22788 44329 22988 44529
rect 23188 44729 23388 44929
rect 22788 44729 22988 44929
rect 16738 49429 16938 49629
rect 17138 49829 17338 50029
rect 23188 45129 23388 45329
rect 22788 45129 22988 45329
rect 23188 45529 23388 45729
rect 22788 45529 22988 45729
rect 23188 45929 23388 46129
rect 22788 45929 22988 46129
rect 23188 46329 23388 46529
rect 22788 46329 22988 46529
rect 23188 33529 23388 33729
rect 22788 33529 22988 33729
rect 23188 33929 23388 34129
rect 22788 33929 22988 34129
rect 23188 34329 23388 34529
rect 22788 34329 22988 34529
rect 23188 34729 23388 34929
rect 22788 34729 22988 34929
rect 23188 35129 23388 35329
rect 22788 35129 22988 35329
rect 23188 35529 23388 35729
rect 22788 35529 22988 35729
rect 23188 35929 23388 36129
rect 22788 35929 22988 36129
rect 23188 36329 23388 36529
rect 22788 36329 22988 36529
rect 23188 36729 23388 36929
rect 22788 36729 22988 36929
rect 23188 37129 23388 37329
rect 22788 37129 22988 37329
rect 23188 37529 23388 37729
rect 22788 37529 22988 37729
rect 23188 37929 23388 38129
rect 22788 37929 22988 38129
rect 23188 38329 23388 38529
rect 22788 38329 22988 38529
rect 23188 38729 23388 38929
rect 22788 38729 22988 38929
rect 23188 39129 23388 39329
rect 22788 39129 22988 39329
rect 23188 39529 23388 39729
rect 22788 39529 22988 39729
rect 23188 39929 23388 40129
rect 22788 39929 22988 40129
rect 23188 40329 23388 40529
rect 22788 40329 22988 40529
rect 23188 40729 23388 40929
rect 22788 40729 22988 40929
rect 23188 41129 23388 41329
rect 22788 41129 22988 41329
rect 23188 41529 23388 41729
rect 22788 41529 22988 41729
rect 23188 28329 23388 28529
rect 22788 28329 22988 28529
rect 23188 28729 23388 28929
rect 22788 28729 22988 28929
rect 23188 29129 23388 29329
rect 22788 29129 22988 29329
rect 23188 29529 23388 29729
rect 22788 29529 22988 29729
rect 23188 29929 23388 30129
rect 22788 29929 22988 30129
rect 23188 30329 23388 30529
rect 22788 30329 22988 30529
rect 23188 30729 23388 30929
rect 22788 30729 22988 30929
rect 23188 31129 23388 31329
rect 22788 31129 22988 31329
rect 23188 31529 23388 31729
rect 22788 31529 22988 31729
rect 23188 31929 23388 32129
rect 22788 31929 22988 32129
rect 23188 32329 23388 32529
rect 22788 32329 22988 32529
rect 23188 32729 23388 32929
rect 22788 32729 22988 32929
rect 23188 33129 23388 33329
rect 22788 33129 22988 33329
rect 44890 17879 45090 18079
rect 44890 17479 45090 17679
rect 47290 17879 47490 18079
rect 47290 17479 47490 17679
rect 46890 17879 47090 18079
rect 46890 17479 47090 17679
rect 46490 17879 46690 18079
rect 46490 17479 46690 17679
rect 46090 17879 46290 18079
rect 46090 17479 46290 17679
rect 45690 17879 45890 18079
rect 45690 17479 45890 17679
rect 45290 17879 45490 18079
rect 45290 17479 45490 17679
rect 47690 17879 47890 18079
rect 47690 17479 47890 17679
rect 32890 17879 33090 18079
rect 32890 17479 33090 17679
rect 32490 17879 32690 18079
rect 32490 17479 32690 17679
rect 32090 17879 32290 18079
rect 32090 17479 32290 17679
rect 31690 17879 31890 18079
rect 31690 17479 31890 17679
rect 31290 17879 31490 18079
rect 31290 17479 31490 17679
rect 30890 17879 31090 18079
rect 44490 17879 44690 18079
rect 44490 17479 44690 17679
rect 44090 17879 44290 18079
rect 44090 17479 44290 17679
rect 43690 17879 43890 18079
rect 43690 17479 43890 17679
rect 43290 17879 43490 18079
rect 43290 17479 43490 17679
rect 42890 17879 43090 18079
rect 42890 17479 43090 17679
rect 42490 17879 42690 18079
rect 42490 17479 42690 17679
rect 42090 17879 42290 18079
rect 42090 17479 42290 17679
rect 41690 17879 41890 18079
rect 41690 17479 41890 17679
rect 41290 17879 41490 18079
rect 41290 17479 41490 17679
rect 40890 17879 41090 18079
rect 40890 17479 41090 17679
rect 40490 17879 40690 18079
rect 40490 17479 40690 17679
rect 40090 17879 40290 18079
rect 40090 17479 40290 17679
rect 39690 17879 39890 18079
rect 39690 17479 39890 17679
rect 39290 17879 39490 18079
rect 39290 17479 39490 17679
rect 38890 17879 39090 18079
rect 38890 17479 39090 17679
rect 38490 17879 38690 18079
rect 38490 17479 38690 17679
rect 38090 17879 38290 18079
rect 38090 17479 38290 17679
rect 37690 17879 37890 18079
rect 37690 17479 37890 17679
rect 37290 17879 37490 18079
rect 37290 17479 37490 17679
rect 36890 17879 37090 18079
rect 36890 17479 37090 17679
rect 36490 17879 36690 18079
rect 36490 17479 36690 17679
rect 36090 17879 36290 18079
rect 36090 17479 36290 17679
rect 35690 17879 35890 18079
rect 35690 17479 35890 17679
rect 35290 17879 35490 18079
rect 35290 17479 35490 17679
rect 34890 17879 35090 18079
rect 34890 17479 35090 17679
rect 34490 17879 34690 18079
rect 34490 17479 34690 17679
rect 34090 17879 34290 18079
rect 34090 17479 34290 17679
rect 33690 17879 33890 18079
rect 33690 17479 33890 17679
rect 33290 17879 33490 18079
rect 33290 17479 33490 17679
rect 30890 17479 31090 17679
rect 30490 17879 30690 18079
rect 30490 17479 30690 17679
rect 30090 17879 30290 18079
rect 30090 17479 30290 17679
rect 23188 14729 23388 14929
rect 22788 14729 22988 14929
rect 23188 15129 23388 15329
rect 22788 15129 22988 15329
rect 23188 15529 23388 15729
rect 22788 15529 22988 15729
rect 22788 24329 22988 24529
rect 23188 24729 23388 24929
rect 23188 15929 23388 16129
rect 22788 15929 22988 16129
rect 23188 16329 23388 16529
rect 22788 16329 22988 16529
rect 23188 16729 23388 16929
rect 22788 16729 22988 16929
rect 23188 17129 23388 17329
rect 22788 17129 22988 17329
rect 23188 17529 23388 17729
rect 22788 17529 22988 17729
rect 23188 17929 23388 18129
rect 22788 17929 22988 18129
rect 23188 18329 23388 18529
rect 22788 18329 22988 18529
rect 23188 18729 23388 18929
rect 22788 18729 22988 18929
rect 23188 19129 23388 19329
rect 22788 19129 22988 19329
rect 23188 26729 23388 26929
rect 22788 26729 22988 26929
rect 23188 27129 23388 27329
rect 22788 27129 22988 27329
rect 23188 27529 23388 27729
rect 22788 27529 22988 27729
rect 23188 19529 23388 19729
rect 23188 24329 23388 24529
rect 27690 17879 27890 18079
rect 27690 17479 27890 17679
rect 27290 17879 27490 18079
rect 27290 17479 27490 17679
rect 26890 17879 27090 18079
rect 26890 17479 27090 17679
rect 26490 17879 26690 18079
rect 26490 17479 26690 17679
rect 26090 17879 26290 18079
rect 26090 17479 26290 17679
rect 25690 17879 25890 18079
rect 25690 17479 25890 17679
rect 25290 17879 25490 18079
rect 25290 17479 25490 17679
rect 22788 26329 22988 26529
rect 23188 23529 23388 23729
rect 22788 23529 22988 23729
rect 23188 23929 23388 24129
rect 22788 23929 22988 24129
rect 22788 23129 22988 23329
rect 23188 14329 23388 14529
rect 22788 14329 22988 14529
rect 29690 17879 29890 18079
rect 29690 17479 29890 17679
rect 29290 17879 29490 18079
rect 29290 17479 29490 17679
rect 28890 17879 29090 18079
rect 28890 17479 29090 17679
rect 28490 17879 28690 18079
rect 28490 17479 28690 17679
rect 28090 17879 28290 18079
rect 28090 17479 28290 17679
rect 22788 24729 22988 24929
rect 23188 25129 23388 25329
rect 22788 25129 22988 25329
rect 23188 25529 23388 25729
rect 22788 25529 22988 25729
rect 23188 25929 23388 26129
rect 22788 25929 22988 26129
rect 23188 26329 23388 26529
rect 22788 19529 22988 19729
rect 23188 19929 23388 20129
rect 22788 19929 22988 20129
rect 23188 20329 23388 20529
rect 22788 20329 22988 20529
rect 23188 20729 23388 20929
rect 22788 20729 22988 20929
rect 23188 21129 23388 21329
rect 22788 21129 22988 21329
rect 23188 21529 23388 21729
rect 22788 21529 22988 21729
rect 23188 21929 23388 22129
rect 22788 21929 22988 22129
rect 23188 22329 23388 22529
rect 22788 22329 22988 22529
rect 23188 22729 23388 22929
rect 22788 22729 22988 22929
rect 23188 23129 23388 23329
rect 23188 8329 23388 8529
rect 22788 8329 22988 8529
rect 23188 8729 23388 8929
rect 22788 8729 22988 8929
rect 23188 9129 23388 9329
rect 22788 9129 22988 9329
rect 23188 9529 23388 9729
rect 22788 9529 22988 9729
rect 23188 9929 23388 10129
rect 22788 9929 22988 10129
rect 23188 10329 23388 10529
rect 22788 10329 22988 10529
rect 23188 10729 23388 10929
rect 22788 10729 22988 10929
rect 23188 11129 23388 11329
rect 22788 11129 22988 11329
rect 23188 11929 23388 12129
rect 22788 11929 22988 12129
rect 23188 12329 23388 12529
rect 22788 12329 22988 12529
rect 23188 12729 23388 12929
rect 22788 12729 22988 12929
rect 23188 13129 23388 13329
rect 22788 13129 22988 13329
rect 23188 13529 23388 13729
rect 22788 13529 22988 13729
rect 23188 13929 23388 14129
rect 22788 13929 22988 14129
rect 23188 7129 23388 7329
rect 22788 7129 22988 7329
rect 23188 7529 23388 7729
rect 22788 7529 22988 7729
rect 23188 7929 23388 8129
rect 22788 7929 22988 8129
rect 23188 11529 23388 11729
rect 22788 11529 22988 11729
rect 66285 27472 66485 27672
rect 66285 27072 66485 27272
rect 69885 27072 70085 27272
rect 69485 27472 69685 27672
rect 69485 27072 69685 27272
rect 69085 27472 69285 27672
rect 69085 27072 69285 27272
rect 68685 27472 68885 27672
rect 68685 27072 68885 27272
rect 68285 27472 68485 27672
rect 68285 27072 68485 27272
rect 67885 27472 68085 27672
rect 67885 27072 68085 27272
rect 67485 27472 67685 27672
rect 67485 27072 67685 27272
rect 67085 27472 67285 27672
rect 67085 27072 67285 27272
rect 66685 27472 66885 27672
rect 66685 27072 66885 27272
rect 70285 27072 70485 27272
rect 69885 27472 70085 27672
rect 73885 27072 74085 27272
rect 73485 27472 73685 27672
rect 73485 27072 73685 27272
rect 73085 27472 73285 27672
rect 73085 27072 73285 27272
rect 72685 27472 72885 27672
rect 72685 27072 72885 27272
rect 72285 27472 72485 27672
rect 72285 27072 72485 27272
rect 71885 27472 72085 27672
rect 71885 27072 72085 27272
rect 71485 27472 71685 27672
rect 71485 27072 71685 27272
rect 71085 27472 71285 27672
rect 71085 27072 71285 27272
rect 70685 27472 70885 27672
rect 83885 27472 84085 27672
rect 83885 27072 84085 27272
rect 83485 27472 83685 27672
rect 83485 27072 83685 27272
rect 83085 27472 83285 27672
rect 83085 27072 83285 27272
rect 82685 27472 82885 27672
rect 82685 27072 82885 27272
rect 82285 27472 82485 27672
rect 82285 27072 82485 27272
rect 81885 27472 82085 27672
rect 81885 27072 82085 27272
rect 81485 27472 81685 27672
rect 81485 27072 81685 27272
rect 81085 27472 81285 27672
rect 81085 27072 81285 27272
rect 80685 27472 80885 27672
rect 80685 27072 80885 27272
rect 80285 27472 80485 27672
rect 80285 27072 80485 27272
rect 79885 27472 80085 27672
rect 79885 27072 80085 27272
rect 79485 27472 79685 27672
rect 79485 27072 79685 27272
rect 79085 27472 79285 27672
rect 79085 27072 79285 27272
rect 78685 27472 78885 27672
rect 78685 27072 78885 27272
rect 78285 27472 78485 27672
rect 78285 27072 78485 27272
rect 77885 27472 78085 27672
rect 77885 27072 78085 27272
rect 77485 27472 77685 27672
rect 77485 27072 77685 27272
rect 77085 27472 77285 27672
rect 77085 27072 77285 27272
rect 76685 27472 76885 27672
rect 76685 27072 76885 27272
rect 76285 27472 76485 27672
rect 76285 27072 76485 27272
rect 75885 27472 76085 27672
rect 75885 27072 76085 27272
rect 75485 27472 75685 27672
rect 75485 27072 75685 27272
rect 75085 27472 75285 27672
rect 75085 27072 75285 27272
rect 74685 27472 74885 27672
rect 74685 27072 74885 27272
rect 74285 27472 74485 27672
rect 74285 27072 74485 27272
rect 73885 27472 74085 27672
rect 70685 27072 70885 27272
rect 70285 27472 70485 27672
rect 52490 17479 52690 17679
rect 52090 17879 52290 18079
rect 54090 17479 54290 17679
rect 65885 27472 66085 27672
rect 65885 27072 66085 27272
rect 65485 27472 65685 27672
rect 65485 27072 65685 27272
rect 53690 17879 53890 18079
rect 53690 17479 53890 17679
rect 53290 17879 53490 18079
rect 53290 17479 53490 17679
rect 52890 17879 53090 18079
rect 48490 17479 48690 17679
rect 64490 17879 64690 18079
rect 64490 17479 64690 17679
rect 64090 17879 64290 18079
rect 64090 17479 64290 17679
rect 63690 17879 63890 18079
rect 63690 17479 63890 17679
rect 63290 17879 63490 18079
rect 63290 17479 63490 17679
rect 62890 17879 63090 18079
rect 62890 17479 63090 17679
rect 62490 17879 62690 18079
rect 62490 17479 62690 17679
rect 62090 17879 62290 18079
rect 62090 17479 62290 17679
rect 61690 17879 61890 18079
rect 61690 17479 61890 17679
rect 61290 17879 61490 18079
rect 61290 17479 61490 17679
rect 60890 17879 61090 18079
rect 60890 17479 61090 17679
rect 60490 17879 60690 18079
rect 60490 17479 60690 17679
rect 52090 17479 52290 17679
rect 52890 17479 53090 17679
rect 52490 17879 52690 18079
rect 51690 17879 51890 18079
rect 51690 17479 51890 17679
rect 51290 17879 51490 18079
rect 51290 17479 51490 17679
rect 50890 17879 51090 18079
rect 50890 17479 51090 17679
rect 50490 17879 50690 18079
rect 50490 17479 50690 17679
rect 50090 17879 50290 18079
rect 50090 17479 50290 17679
rect 49690 17879 49890 18079
rect 49690 17479 49890 17679
rect 49290 17879 49490 18079
rect 49290 17479 49490 17679
rect 48890 17879 49090 18079
rect 48890 17479 49090 17679
rect 48490 17879 48690 18079
rect 60090 17879 60290 18079
rect 60090 17479 60290 17679
rect 59690 17879 59890 18079
rect 59690 17479 59890 17679
rect 59290 17879 59490 18079
rect 59290 17479 59490 17679
rect 58890 17879 59090 18079
rect 58890 17479 59090 17679
rect 58490 17879 58690 18079
rect 58490 17479 58690 17679
rect 58090 17879 58290 18079
rect 58090 17479 58290 17679
rect 57690 17879 57890 18079
rect 57690 17479 57890 17679
rect 57290 17879 57490 18079
rect 57290 17479 57490 17679
rect 56890 17879 57090 18079
rect 56890 17479 57090 17679
rect 56490 17879 56690 18079
rect 56490 17479 56690 17679
rect 56090 17879 56290 18079
rect 56090 17479 56290 17679
rect 55690 17879 55890 18079
rect 55690 17479 55890 17679
rect 55290 17879 55490 18079
rect 55290 17479 55490 17679
rect 54890 17879 55090 18079
rect 54890 17479 55090 17679
rect 54490 17879 54690 18079
rect 54490 17479 54690 17679
rect 54090 17879 54290 18079
rect 156820 27860 157020 28060
rect 156020 27860 156220 28060
rect 155620 27860 155820 28060
rect 156420 27860 156620 28060
rect 156020 41860 156220 42060
rect 155620 41860 155820 42060
rect 156420 41860 156620 42060
rect 156820 41860 157020 42060
rect 156020 48660 156220 48860
rect 156420 48660 156620 48860
rect 155620 48660 155820 48860
rect 156820 48660 157020 48860
rect 156420 50260 156620 50460
rect 156020 54660 156220 54860
rect 156420 51060 156620 51260
rect 156420 49860 156620 50060
rect 156020 52660 156220 52860
rect 156420 49460 156620 49660
rect 156420 49060 156620 49260
rect 156420 50660 156620 50860
rect 156020 52260 156220 52460
rect 156020 54260 156220 54460
rect 155620 55460 155820 55660
rect 156020 51860 156220 52060
rect 155620 55060 155820 55260
rect 156420 55460 156620 55660
rect 155620 54660 155820 54860
rect 156420 55060 156620 55260
rect 156820 55460 157020 55660
rect 155620 54260 155820 54460
rect 156820 55060 157020 55260
rect 155620 53860 155820 54060
rect 156020 51460 156220 51660
rect 156420 54660 156620 54860
rect 156820 54660 157020 54860
rect 155620 53460 155820 53660
rect 156420 54260 156620 54460
rect 156820 54260 157020 54460
rect 155620 53060 155820 53260
rect 156820 53860 157020 54060
rect 155620 52660 155820 52860
rect 156020 51060 156220 51260
rect 156420 53860 156620 54060
rect 156820 53460 157020 53660
rect 156020 53860 156220 54060
rect 155620 52260 155820 52460
rect 156420 53460 156620 53660
rect 156820 53060 157020 53260
rect 155620 51860 155820 52060
rect 156820 52660 157020 52860
rect 155620 51460 155820 51660
rect 156020 55060 156220 55260
rect 156420 53060 156620 53260
rect 156020 50660 156220 50860
rect 156820 52260 157020 52460
rect 155620 51060 155820 51260
rect 156820 51860 157020 52060
rect 156420 52660 156620 52860
rect 155620 50660 155820 50860
rect 156820 51460 157020 51660
rect 155620 50260 155820 50460
rect 156820 51060 157020 51260
rect 155620 49860 155820 50060
rect 156420 52260 156620 52460
rect 156820 50660 157020 50860
rect 155620 49460 155820 49660
rect 156020 50260 156220 50460
rect 156820 50260 157020 50460
rect 155620 49060 155820 49260
rect 156020 53460 156220 53660
rect 156020 49460 156220 49660
rect 156820 49860 157020 50060
rect 156420 51860 156620 52060
rect 156020 55460 156220 55660
rect 156820 49460 157020 49660
rect 156020 49860 156220 50060
rect 156820 49060 157020 49260
rect 156420 51460 156620 51660
rect 156020 49060 156220 49260
rect 156020 53060 156220 53260
rect 156420 47060 156620 47260
rect 156820 47460 157020 47660
rect 156820 46660 157020 46860
rect 156020 44660 156220 44860
rect 156420 44260 156620 44460
rect 156020 46260 156220 46460
rect 156820 43860 157020 44060
rect 156020 42260 156220 42460
rect 156420 46660 156620 46860
rect 156820 43060 157020 43260
rect 156420 43860 156620 44060
rect 155620 44260 155820 44460
rect 156020 44260 156220 44460
rect 156820 45060 157020 45260
rect 156820 47860 157020 48060
rect 156020 47460 156220 47660
rect 155620 46260 155820 46460
rect 155620 42660 155820 42860
rect 156420 43460 156620 43660
rect 156420 48260 156620 48460
rect 156420 46260 156620 46460
rect 155620 46660 155820 46860
rect 156020 43860 156220 44060
rect 156420 43060 156620 43260
rect 156020 45860 156220 46060
rect 155620 45460 155820 45660
rect 156820 44260 157020 44460
rect 156820 45860 157020 46060
rect 156420 42660 156620 42860
rect 156020 47060 156220 47260
rect 156820 42660 157020 42860
rect 156420 47860 156620 48060
rect 156420 42260 156620 42460
rect 156020 43460 156220 43660
rect 156420 45860 156620 46060
rect 156820 46260 157020 46460
rect 155620 43860 155820 44060
rect 155620 45860 155820 46060
rect 155620 43060 155820 43260
rect 156020 45460 156220 45660
rect 156420 45460 156620 45660
rect 155620 44660 155820 44860
rect 156820 44660 157020 44860
rect 156420 47460 156620 47660
rect 156020 43060 156220 43260
rect 156820 43460 157020 43660
rect 156020 47860 156220 48060
rect 156820 42260 157020 42460
rect 155620 45060 155820 45260
rect 155620 42260 155820 42460
rect 156420 45060 156620 45260
rect 156020 45060 156220 45260
rect 155620 48260 155820 48460
rect 156020 46660 156220 46860
rect 155620 43460 155820 43660
rect 156020 42660 156220 42860
rect 155620 47860 155820 48060
rect 156020 48260 156220 48460
rect 155620 47060 155820 47260
rect 155620 47460 155820 47660
rect 156820 47060 157020 47260
rect 156420 44660 156620 44860
rect 156820 45460 157020 45660
rect 156820 48260 157020 48460
rect 156020 35060 156220 35260
rect 155620 36660 155820 36860
rect 156820 41460 157020 41660
rect 156420 39460 156620 39660
rect 155620 35460 155820 35660
rect 156820 41060 157020 41260
rect 155620 40660 155820 40860
rect 155620 39460 155820 39660
rect 156820 38260 157020 38460
rect 156020 40660 156220 40860
rect 156420 40660 156620 40860
rect 156420 37060 156620 37260
rect 156020 38260 156220 38460
rect 155620 41060 155820 41260
rect 155620 37060 155820 37260
rect 156820 36260 157020 36460
rect 156020 39860 156220 40060
rect 155620 35060 155820 35260
rect 156820 35060 157020 35260
rect 156420 39060 156620 39260
rect 156820 39860 157020 40060
rect 156420 35060 156620 35260
rect 156420 41060 156620 41260
rect 156420 40260 156620 40460
rect 156820 38660 157020 38860
rect 156420 41460 156620 41660
rect 156420 37860 156620 38060
rect 156020 37060 156220 37260
rect 155620 37460 155820 37660
rect 156020 37460 156220 37660
rect 156820 37860 157020 38060
rect 156020 41460 156220 41660
rect 156820 35860 157020 36060
rect 156420 36660 156620 36860
rect 156420 35860 156620 36060
rect 156020 37860 156220 38060
rect 155620 39860 155820 40060
rect 155620 40260 155820 40460
rect 156420 37460 156620 37660
rect 156820 36660 157020 36860
rect 156420 39860 156620 40060
rect 155620 41460 155820 41660
rect 156020 36660 156220 36860
rect 156420 38660 156620 38860
rect 155620 38660 155820 38860
rect 156020 39460 156220 39660
rect 156820 37460 157020 37660
rect 156020 36260 156220 36460
rect 156820 40260 157020 40460
rect 156420 35460 156620 35660
rect 155620 36260 155820 36460
rect 156820 39460 157020 39660
rect 156020 40260 156220 40460
rect 155620 38260 155820 38460
rect 156020 41060 156220 41260
rect 156020 35860 156220 36060
rect 156420 38260 156620 38460
rect 156020 39060 156220 39260
rect 156820 37060 157020 37260
rect 155620 35860 155820 36060
rect 156020 35460 156220 35660
rect 155620 39060 155820 39260
rect 156820 40660 157020 40860
rect 156420 36260 156620 36460
rect 156820 39060 157020 39260
rect 156820 35460 157020 35660
rect 156020 38660 156220 38860
rect 155620 37860 155820 38060
rect 156020 33860 156220 34060
rect 156420 33460 156620 33660
rect 155620 31460 155820 31660
rect 156820 29060 157020 29260
rect 156820 31060 157020 31260
rect 155620 28660 155820 28860
rect 156820 33060 157020 33260
rect 156020 31060 156220 31260
rect 155620 34660 155820 34860
rect 156020 32260 156220 32460
rect 156420 34660 156620 34860
rect 156420 29460 156620 29660
rect 156420 33860 156620 34060
rect 156420 30260 156620 30460
rect 156820 28660 157020 28860
rect 156020 33460 156220 33660
rect 156820 33860 157020 34060
rect 156420 28260 156620 28460
rect 155620 32660 155820 32860
rect 156420 31460 156620 31660
rect 156420 32660 156620 32860
rect 156420 30660 156620 30860
rect 156420 29860 156620 30060
rect 156020 28660 156220 28860
rect 156420 28660 156620 28860
rect 155620 31860 155820 32060
rect 156020 34660 156220 34860
rect 155620 29060 155820 29260
rect 155620 30260 155820 30460
rect 155620 33060 155820 33260
rect 156420 34260 156620 34460
rect 156420 31060 156620 31260
rect 156020 34260 156220 34460
rect 156420 33060 156620 33260
rect 156820 33460 157020 33660
rect 155620 31060 155820 31260
rect 156020 33060 156220 33260
rect 156020 31460 156220 31660
rect 156820 34260 157020 34460
rect 156820 30660 157020 30860
rect 156820 34660 157020 34860
rect 156020 32660 156220 32860
rect 156020 28260 156220 28460
rect 156820 29860 157020 30060
rect 156820 28260 157020 28460
rect 155620 33460 155820 33660
rect 155620 30660 155820 30860
rect 156820 32260 157020 32460
rect 156020 31860 156220 32060
rect 156020 29060 156220 29260
rect 156420 29060 156620 29260
rect 155620 34260 155820 34460
rect 156420 31860 156620 32060
rect 156020 30260 156220 30460
rect 156020 30660 156220 30860
rect 155620 29860 155820 30060
rect 156820 31460 157020 31660
rect 156820 29460 157020 29660
rect 156420 32260 156620 32460
rect 156020 29460 156220 29660
rect 155620 33860 155820 34060
rect 155620 28260 155820 28460
rect 155620 32260 155820 32460
rect 156820 31860 157020 32060
rect 155620 29460 155820 29660
rect 156820 30260 157020 30460
rect 156020 29860 156220 30060
rect 156820 32660 157020 32860
rect 99415 49559 99615 49759
rect 99415 50759 99615 50959
rect 99815 53159 100015 53359
rect 99815 51159 100015 51359
rect 99415 53159 99615 53359
rect 99815 53559 100015 53759
rect 99815 49959 100015 50159
rect 99415 53559 99615 53759
rect 99815 54359 100015 54559
rect 99415 54359 99615 54559
rect 99815 54759 100015 54959
rect 99415 51159 99615 51359
rect 99415 54759 99615 54959
rect 99815 51559 100015 51759
rect 99415 55559 99615 55759
rect 99815 55159 100015 55359
rect 99415 51559 99615 51759
rect 99415 49959 99615 50159
rect 99815 50359 100015 50559
rect 99815 51959 100015 52159
rect 99815 53959 100015 54159
rect 99415 55159 99615 55359
rect 99815 55559 100015 55759
rect 99415 51959 99615 52159
rect 99815 52359 100015 52559
rect 99415 50359 99615 50559
rect 99815 49559 100015 49759
rect 99415 53959 99615 54159
rect 99415 52359 99615 52559
rect 99815 52759 100015 52959
rect 99815 50759 100015 50959
rect 99415 52759 99615 52959
rect 103485 27072 103685 27272
rect 103085 27472 103285 27672
rect 103085 27072 103285 27272
rect 102685 27472 102885 27672
rect 102685 27072 102885 27272
rect 104685 27472 104885 27672
rect 104685 27072 104885 27272
rect 104285 27472 104485 27672
rect 104285 27072 104485 27272
rect 103885 27472 104085 27672
rect 103885 27072 104085 27272
rect 103485 27472 103685 27672
rect 85085 27072 85285 27272
rect 100285 27472 100485 27672
rect 91885 27072 92085 27272
rect 93885 27072 94085 27272
rect 99885 27072 100085 27272
rect 99485 27472 99685 27672
rect 93485 27472 93685 27672
rect 85485 27472 85685 27672
rect 88685 27472 88885 27672
rect 102285 27472 102485 27672
rect 91485 27472 91685 27672
rect 99485 27072 99685 27272
rect 91485 27072 91685 27272
rect 85485 27072 85685 27272
rect 99085 27472 99285 27672
rect 93085 27072 93285 27272
rect 92685 27472 92885 27672
rect 102285 27072 102485 27272
rect 101885 27472 102085 27672
rect 91085 27472 91285 27672
rect 99085 27072 99285 27272
rect 98685 27472 98885 27672
rect 91085 27072 91285 27272
rect 94685 27072 94885 27272
rect 101885 27072 102085 27272
rect 88285 27472 88485 27672
rect 88285 27072 88485 27272
rect 98685 27072 98885 27272
rect 98285 27472 98485 27672
rect 101485 27472 101685 27672
rect 90685 27472 90885 27672
rect 87085 27472 87285 27672
rect 101485 27072 101685 27272
rect 90685 27072 90885 27272
rect 98285 27072 98485 27272
rect 101085 27472 101285 27672
rect 87085 27072 87285 27272
rect 97885 27472 98085 27672
rect 94285 27072 94485 27272
rect 87885 27472 88085 27672
rect 101085 27072 101285 27272
rect 90285 27472 90485 27672
rect 84685 27472 84885 27672
rect 97885 27072 98085 27272
rect 97485 27472 97685 27672
rect 100685 27472 100885 27672
rect 87885 27072 88085 27272
rect 100685 27072 100885 27272
rect 93885 27472 94085 27672
rect 94285 27472 94485 27672
rect 97485 27072 97685 27272
rect 97085 27472 97285 27672
rect 84685 27072 84885 27272
rect 90285 27072 90485 27272
rect 92285 27072 92485 27272
rect 95485 27072 95685 27272
rect 88685 27072 88885 27272
rect 97085 27072 97285 27272
rect 85085 27472 85285 27672
rect 92685 27072 92885 27272
rect 96685 27472 96885 27672
rect 89885 27472 90085 27672
rect 86685 27472 86885 27672
rect 86685 27072 86885 27272
rect 89885 27072 90085 27272
rect 85885 27472 86085 27672
rect 96685 27072 96885 27272
rect 96285 27472 96485 27672
rect 85885 27072 86085 27272
rect 92285 27472 92485 27672
rect 93485 27072 93685 27272
rect 93085 27472 93285 27672
rect 89485 27472 89685 27672
rect 96285 27072 96485 27272
rect 95885 27472 96085 27672
rect 89485 27072 89685 27272
rect 87485 27072 87685 27272
rect 100285 27072 100485 27272
rect 95085 27072 95285 27272
rect 86285 27472 86485 27672
rect 86285 27072 86485 27272
rect 89085 27472 89285 27672
rect 89085 27072 89285 27272
rect 95885 27072 96085 27272
rect 99885 27472 100085 27672
rect 95485 27472 95685 27672
rect 91885 27472 92085 27672
rect 94685 27472 94885 27672
rect 95085 27472 95285 27672
rect 87485 27472 87685 27672
rect 156420 21060 156620 21260
rect 156820 21060 157020 21260
rect 156020 21060 156220 21260
rect 155620 21060 155820 21260
rect 156020 25460 156220 25660
rect 156020 23860 156220 24060
rect 155620 24660 155820 24860
rect 156420 23060 156620 23260
rect 156420 22260 156620 22460
rect 156020 22260 156220 22460
rect 155620 26660 155820 26860
rect 156820 27460 157020 27660
rect 155620 24260 155820 24460
rect 156020 27060 156220 27260
rect 156820 22660 157020 22860
rect 156020 27460 156220 27660
rect 156020 22660 156220 22860
rect 156420 26660 156620 26860
rect 155620 23860 155820 24060
rect 156820 23460 157020 23660
rect 156820 27060 157020 27260
rect 156020 23060 156220 23260
rect 156020 21460 156220 21660
rect 155620 26260 155820 26460
rect 156420 23860 156620 24060
rect 156020 24660 156220 24860
rect 156820 25060 157020 25260
rect 156820 22260 157020 22460
rect 155620 23460 155820 23660
rect 155620 25060 155820 25260
rect 155620 21460 155820 21660
rect 156820 26660 157020 26860
rect 156420 21860 156620 22060
rect 156420 23460 156620 23660
rect 155620 23060 155820 23260
rect 156820 26260 157020 26460
rect 156420 27060 156620 27260
rect 156020 26260 156220 26460
rect 156420 26260 156620 26460
rect 156020 23460 156220 23660
rect 155620 25860 155820 26060
rect 155620 22660 155820 22860
rect 156420 24660 156620 24860
rect 156820 21860 157020 22060
rect 156020 26660 156220 26860
rect 156020 25860 156220 26060
rect 156420 27460 156620 27660
rect 156020 24260 156220 24460
rect 155620 27460 155820 27660
rect 156820 25860 157020 26060
rect 156420 22660 156620 22860
rect 155620 22260 155820 22460
rect 156020 25060 156220 25260
rect 156020 21860 156220 22060
rect 156820 21460 157020 21660
rect 156820 23060 157020 23260
rect 156420 25460 156620 25660
rect 155620 21860 155820 22060
rect 156820 25460 157020 25660
rect 156420 25060 156620 25260
rect 156420 21460 156620 21660
rect 156820 23860 157020 24060
rect 156420 24260 156620 24460
rect 156820 24260 157020 24460
rect 156420 25860 156620 26060
rect 155620 25460 155820 25660
rect 155620 27060 155820 27260
rect 156820 24660 157020 24860
rect 156020 18660 156220 18860
rect 155620 18660 155820 18860
rect 156420 14260 156620 14460
rect 156020 20260 156220 20460
rect 156420 15860 156620 16060
rect 156820 18260 157020 18460
rect 155620 17860 155820 18060
rect 156420 20660 156620 20860
rect 156820 17060 157020 17260
rect 156020 19860 156220 20060
rect 155620 19460 155820 19660
rect 156020 14260 156220 14460
rect 155620 18260 155820 18460
rect 156820 15060 157020 15260
rect 156820 14660 157020 14860
rect 155620 16260 155820 16460
rect 155620 15460 155820 15660
rect 156020 19460 156220 19660
rect 155620 17060 155820 17260
rect 156020 16660 156220 16860
rect 156820 19860 157020 20060
rect 156020 19060 156220 19260
rect 156420 19460 156620 19660
rect 155620 19060 155820 19260
rect 156020 17860 156220 18060
rect 156820 19460 157020 19660
rect 156420 17060 156620 17260
rect 156820 16660 157020 16860
rect 156020 18260 156220 18460
rect 156820 20660 157020 20860
rect 156420 18660 156620 18860
rect 156820 15460 157020 15660
rect 156020 15460 156220 15660
rect 156420 16260 156620 16460
rect 156420 17860 156620 18060
rect 156820 20260 157020 20460
rect 156020 15060 156220 15260
rect 156420 20260 156620 20460
rect 156420 15460 156620 15660
rect 155620 17460 155820 17660
rect 156420 18260 156620 18460
rect 156420 16660 156620 16860
rect 156820 19060 157020 19260
rect 156820 15860 157020 16060
rect 156420 15060 156620 15260
rect 156820 16260 157020 16460
rect 156020 16260 156220 16460
rect 156820 17460 157020 17660
rect 155620 15860 155820 16060
rect 156420 19060 156620 19260
rect 155620 14660 155820 14860
rect 156020 17060 156220 17260
rect 155620 20660 155820 20860
rect 156020 17460 156220 17660
rect 156020 15860 156220 16060
rect 156820 18660 157020 18860
rect 156020 14660 156220 14860
rect 156420 19860 156620 20060
rect 155620 15060 155820 15260
rect 155620 20260 155820 20460
rect 156820 17860 157020 18060
rect 156820 14260 157020 14460
rect 155620 19860 155820 20060
rect 155620 14260 155820 14460
rect 156420 14660 156620 14860
rect 156020 20660 156220 20860
rect 156420 17460 156620 17660
rect 155620 16660 155820 16860
rect 156820 7060 157020 7260
rect 156420 7060 156620 7260
rect 155620 7060 155820 7260
rect 156020 7060 156220 7260
rect 156020 10660 156220 10860
rect 156420 8660 156620 8860
rect 156820 12660 157020 12860
rect 155620 12260 155820 12460
rect 156820 13460 157020 13660
rect 156020 7860 156220 8060
rect 155620 11460 155820 11660
rect 155620 10260 155820 10460
rect 156820 11060 157020 11260
rect 155620 9060 155820 9260
rect 156820 7460 157020 7660
rect 156020 13060 156220 13260
rect 156020 8260 156220 8460
rect 155620 10660 155820 10860
rect 156020 12660 156220 12860
rect 156420 10660 156620 10860
rect 156020 9460 156220 9660
rect 156820 11460 157020 11660
rect 156820 13860 157020 14060
rect 155620 13860 155820 14060
rect 156420 8260 156620 8460
rect 156420 9860 156620 10060
rect 156020 11860 156220 12060
rect 156820 10260 157020 10460
rect 156020 9860 156220 10060
rect 156420 9060 156620 9260
rect 156420 11460 156620 11660
rect 156820 9860 157020 10060
rect 156420 13060 156620 13260
rect 155620 12660 155820 12860
rect 155620 9860 155820 10060
rect 156420 10260 156620 10460
rect 156820 9060 157020 9260
rect 155620 11860 155820 12060
rect 156020 7460 156220 7660
rect 156020 13460 156220 13660
rect 156020 11060 156220 11260
rect 156420 13460 156620 13660
rect 156420 12260 156620 12460
rect 155620 13460 155820 13660
rect 156820 7860 157020 8060
rect 156820 9460 157020 9660
rect 156420 13860 156620 14060
rect 155620 7860 155820 8060
rect 156020 9060 156220 9260
rect 155620 8260 155820 8460
rect 156020 13860 156220 14060
rect 156420 11860 156620 12060
rect 156820 13060 157020 13260
rect 156820 10660 157020 10860
rect 155620 13060 155820 13260
rect 156020 8660 156220 8860
rect 156820 8260 157020 8460
rect 155620 8660 155820 8860
rect 156420 11060 156620 11260
rect 156020 10260 156220 10460
rect 156420 9460 156620 9660
rect 156420 12660 156620 12860
rect 156420 7460 156620 7660
rect 156020 12260 156220 12460
rect 156820 12260 157020 12460
rect 156820 8660 157020 8860
rect 155620 7460 155820 7660
rect 156820 11860 157020 12060
rect 155620 11060 155820 11260
rect 156020 11460 156220 11660
rect 155620 9460 155820 9660
rect 156420 7860 156620 8060
rect 155620 2260 155820 2460
rect 156020 2660 156220 2860
rect 156420 3460 156620 3660
rect 156420 4660 156620 4860
rect 155620 4260 155820 4460
rect 155620 1060 155820 1260
rect 156020 4660 156220 4860
rect 156420 5460 156620 5660
rect 156420 2260 156620 2460
rect 155620 2660 155820 2860
rect 156820 1460 157020 1660
rect 156820 5060 157020 5260
rect 156820 2660 157020 2860
rect 156820 1860 157020 2060
rect 156020 5860 156220 6060
rect 156420 3060 156620 3260
rect 155620 5060 155820 5260
rect 155620 660 155820 860
rect 156820 660 157020 860
rect 156820 1060 157020 1260
rect 156020 3060 156220 3260
rect 156420 1060 156620 1260
rect 156420 6660 156620 6860
rect 156820 5460 157020 5660
rect 156020 6260 156220 6460
rect 155620 6660 155820 6860
rect 156420 6260 156620 6460
rect 155620 3460 155820 3660
rect 155620 3060 155820 3260
rect 156420 5860 156620 6060
rect 156820 3060 157020 3260
rect 155620 6260 155820 6460
rect 155620 260 155820 460
rect 156020 2260 156220 2460
rect 156820 4660 157020 4860
rect 156420 1860 156620 2060
rect 156420 260 156620 460
rect 155620 1860 155820 2060
rect 156020 6660 156220 6860
rect 156020 3460 156220 3660
rect 156420 2660 156620 2860
rect 156020 1860 156220 2060
rect 156020 260 156220 460
rect 155620 3860 155820 4060
rect 156420 3860 156620 4060
rect 156820 2260 157020 2460
rect 156820 3460 157020 3660
rect 155620 4660 155820 4860
rect 156420 660 156620 860
rect 155620 1460 155820 1660
rect 156820 6260 157020 6460
rect 156020 1060 156220 1260
rect 156020 5060 156220 5260
rect 156820 4260 157020 4460
rect 156820 3860 157020 4060
rect 156420 4260 156620 4460
rect 156020 660 156220 860
rect 156820 6660 157020 6860
rect 156020 4260 156220 4460
rect 156020 3860 156220 4060
rect 156820 5860 157020 6060
rect 156420 1460 156620 1660
rect 156020 5460 156220 5660
rect 156820 260 157020 460
rect 155620 5860 155820 6060
rect 155620 5460 155820 5660
rect 156020 1460 156220 1660
rect 156420 5060 156620 5260
<< l71d20 >>
rect 0 0 2000 111520
rect 155320 0 157320 111520
<< l70d20 >>
rect 21430 106848 41130 111520
rect 107186 101982 109356 102352
rect 0 0 153165 106848
rect 0 106848 21430 111520
rect 139578 106848 153165 111520
rect 155320 0 157320 111520
<< l71d16 >>
rect 155320 0 157320 111520
rect 134630 110520 134930 111520
rect 137390 110520 137690 111520
rect 131870 110520 132170 111520
rect 129110 110520 129410 111520
rect 126350 110520 126650 111520
rect 123590 110520 123890 111520
rect 120830 110520 121130 111520
rect 118070 110520 118370 111520
rect 115310 110520 115610 111520
rect 112550 110520 112850 111520
rect 109790 110520 110090 111520
rect 107030 110520 107330 111520
rect 104270 110520 104570 111520
rect 101510 110520 101810 111520
rect 98750 110520 99050 111520
rect 95990 110520 96290 111520
rect 93230 110520 93530 111520
rect 90470 110520 90770 111520
rect 87710 110520 88010 111520
rect 40790 110520 41090 111520
rect 38030 110520 38330 111520
rect 35270 110520 35570 111520
rect 32510 110520 32810 111520
rect 29750 110520 30050 111520
rect 26990 110520 27290 111520
rect 24230 110520 24530 111520
rect 21470 110520 21770 111520
rect 62870 110520 63170 111520
rect 60110 110520 60410 111520
rect 57350 110520 57650 111520
rect 54590 110520 54890 111520
rect 51830 110520 52130 111520
rect 49070 110520 49370 111520
rect 46310 110520 46610 111520
rect 43550 110520 43850 111520
rect 84950 110520 85250 111520
rect 82190 110520 82490 111520
rect 79430 110520 79730 111520
rect 76670 110520 76970 111520
rect 0 0 2000 111520
rect 73910 110520 74210 111520
rect 71150 110520 71450 111520
rect 68390 110520 68690 111520
rect 65630 110520 65930 111520
<< labels >>
rlabel l71d5 156337 58314 156337 58314 0 VGND
rlabel l71d5 134780 111020 134780 111020 0 clk
rlabel l71d5 137540 111020 137540 111020 0 ena
rlabel l71d5 132020 111020 132020 111020 0 rst_n
rlabel l71d5 129260 111020 129260 111020 0 ui_in[0]
rlabel l71d5 126500 111020 126500 111020 0 ui_in[1]
rlabel l71d5 123740 111020 123740 111020 0 ui_in[2]
rlabel l71d5 120980 111020 120980 111020 0 ui_in[3]
rlabel l71d5 118220 111020 118220 111020 0 ui_in[4]
rlabel l71d5 115460 111020 115460 111020 0 ui_in[5]
rlabel l71d5 112700 111020 112700 111020 0 ui_in[6]
rlabel l71d5 109940 111020 109940 111020 0 ui_in[7]
rlabel l71d5 107180 111020 107180 111020 0 uio_in[0]
rlabel l71d5 104420 111020 104420 111020 0 uio_in[1]
rlabel l71d5 101660 111020 101660 111020 0 uio_in[2]
rlabel l71d5 98900 111020 98900 111020 0 uio_in[3]
rlabel l71d5 96140 111020 96140 111020 0 uio_in[4]
rlabel l71d5 93380 111020 93380 111020 0 uio_in[5]
rlabel l71d5 90620 111020 90620 111020 0 uio_in[6]
rlabel l71d5 87860 111020 87860 111020 0 uio_in[7]
rlabel l71d5 40940 111020 40940 111020 0 uio_oe[0]
rlabel l71d5 38180 111020 38180 111020 0 uio_oe[1]
rlabel l71d5 35420 111020 35420 111020 0 uio_oe[2]
rlabel l71d5 32660 111020 32660 111020 0 uio_oe[3]
rlabel l71d5 29900 111020 29900 111020 0 uio_oe[4]
rlabel l71d5 27140 111020 27140 111020 0 uio_oe[5]
rlabel l71d5 24380 111020 24380 111020 0 uio_oe[6]
rlabel l71d5 21620 111020 21620 111020 0 uio_oe[7]
rlabel l71d5 63020 111020 63020 111020 0 uio_out[0]
rlabel l71d5 60260 111020 60260 111020 0 uio_out[1]
rlabel l71d5 57500 111020 57500 111020 0 uio_out[2]
rlabel l71d5 54740 111020 54740 111020 0 uio_out[3]
rlabel l71d5 51980 111020 51980 111020 0 uio_out[4]
rlabel l71d5 49220 111020 49220 111020 0 uio_out[5]
rlabel l71d5 46460 111020 46460 111020 0 uio_out[6]
rlabel l71d5 43700 111020 43700 111020 0 uio_out[7]
rlabel l71d5 85100 111020 85100 111020 0 uo_out[0]
rlabel l71d5 82340 111020 82340 111020 0 uo_out[1]
rlabel l71d5 79580 111020 79580 111020 0 uo_out[2]
rlabel l71d5 76820 111020 76820 111020 0 uo_out[3]
rlabel l71d5 74060 111020 74060 111020 0 uo_out[4]
rlabel l71d5 71300 111020 71300 111020 0 uo_out[5]
rlabel l71d5 68540 111020 68540 111020 0 uo_out[6]
rlabel l71d5 65780 111020 65780 111020 0 uo_out[7]
rlabel l71d5 1114 60965 1114 60965 0 VPWR
use dac_8bit dac_8bit_1
timestamp 1698899266
transform 0 -1 132001 -1 0 107532
box -350 -90 7270 25260
use inv_strvd inv_strvd_1
timestamp 1698899266
transform -1 0 85420 0 1 16174
box -20590 -789 20615 12166
use driver driver_1
timestamp 1698899266
transform -1 0 308467 0 -1 306887
box 205776 200205 223200 203405
use inv_strvd inv_strvd_2
timestamp 1698899266
transform 0 1 5840 1 0 67694
box -20590 -789 20615 12166
use inv_strvd inv_strvd_3
timestamp 1698899266
transform 0 -1 110913 -1 0 69494
box -20590 -789 20615 12166
use inv_strvd inv_strvd_4
timestamp 1698899266
transform -1 0 45225 0 1 6581
box -20590 -789 20615 12166
use inv_strvd inv_strvd_5
timestamp 1698899266
transform 1 0 76545 0 -1 100625
box -20590 -789 20615 12166
use inv_strvd inv_strvd_6
timestamp 1698899266
transform 1 0 31335 0 -1 102525
box -20590 -789 20615 12166
use inv_strvd inv_strvd_7
timestamp 1698899266
transform 0 1 11890 1 0 26594
box -20590 -789 20615 12166
use pin_connect pin_connect_1
timestamp 1698899266
transform 1 0 21435 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_2
timestamp 1698899266
transform 1 0 24195 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_3
timestamp 1698899266
transform 1 0 26955 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_4
timestamp 1698899266
transform 1 0 29715 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_5
timestamp 1698899266
transform 1 0 32475 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_6
timestamp 1698899266
transform 1 0 35235 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_7
timestamp 1698899266
transform 1 0 37995 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_8
timestamp 1698899266
transform 1 0 40755 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_9
timestamp 1698899266
transform 1 0 43515 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_10
timestamp 1698899266
transform 1 0 46275 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_11
timestamp 1698899266
transform 1 0 49035 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_12
timestamp 1698899266
transform 1 0 51795 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_13
timestamp 1698899266
transform 1 0 54555 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_14
timestamp 1698899266
transform 1 0 57315 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_15
timestamp 1698899266
transform 1 0 60075 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_16
timestamp 1698899266
transform 1 0 62835 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_17
timestamp 1698899266
transform 1 0 65595 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_18
timestamp 1698899266
transform 1 0 68355 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_19
timestamp 1698899266
transform 1 0 71115 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_20
timestamp 1698899266
transform 1 0 73875 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_21
timestamp 1698899266
transform 1 0 76635 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_22
timestamp 1698899266
transform 1 0 79395 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_23
timestamp 1698899266
transform 1 0 82155 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_24
timestamp 1698899266
transform 1 0 84915 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_25
timestamp 1698899266
transform 1 0 87675 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_26
timestamp 1698899266
transform 1 0 90435 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_27
timestamp 1698899266
transform 1 0 93195 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_28
timestamp 1698899266
transform 1 0 95955 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_29
timestamp 1698899266
transform 1 0 98715 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_30
timestamp 1698899266
transform 1 0 101475 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_31
timestamp 1698899266
transform 1 0 104235 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_32
timestamp 1698899266
transform 1 0 106995 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_33
timestamp 1698899266
transform 1 0 109755 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_34
timestamp 1698899266
transform 1 0 112515 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_35
timestamp 1698899266
transform 1 0 115275 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_36
timestamp 1698899266
transform 1 0 118035 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_37
timestamp 1698899266
transform 1 0 120795 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_38
timestamp 1698899266
transform 1 0 123555 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_39
timestamp 1698899266
transform 1 0 126315 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_40
timestamp 1698899266
transform 1 0 129075 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_41
timestamp 1698899266
transform 1 0 131835 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_42
timestamp 1698899266
transform 1 0 134595 0 1 108928
box -5 0 375 2592
use pin_connect pin_connect_43
timestamp 1698899266
transform 1 0 137355 0 1 108928
box -5 0 375 2592
use tt_um_template tt_um_template_1
timestamp 1698899266
transform 1 0 0 0 1 0
box 0 0 157320 111520
<< end >>
