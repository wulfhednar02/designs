magic
tech sky130A
timestamp 1698982078
<< end >>
