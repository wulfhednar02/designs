magic
tech sky130A
magscale 1 2
timestamp 1699066547
<< error_s >>
rect 17141 21212 17153 21218
rect 17163 21194 17165 21206
rect 20416 21122 20422 21128
rect 20386 21098 20392 21118
rect 20344 21010 20350 21030
rect 20386 20988 20392 20994
rect 17163 20826 17165 20838
rect 17141 20814 17153 20820
rect 2298 20388 2498 20410
rect 21916 20398 21944 20468
rect 22910 20398 22938 20468
rect 23904 20398 23932 20468
rect 24898 20398 24926 20468
rect 22413 20144 22441 20214
rect 23407 20144 23435 20214
rect 24401 20144 24429 20214
rect 25395 20144 25423 20214
rect 11340 20008 11540 20030
rect 2288 19666 8340 19667
rect 11330 19286 17382 19287
rect 21302 17852 21345 17920
rect 1317 9586 1339 9824
rect 2006 9586 2049 15654
rect 21344 11826 21345 17852
rect 22066 17668 22088 17868
rect 2006 9560 2007 9586
rect 2527 1366 2549 1604
rect 3216 1366 3259 7434
rect 14969 4073 21105 4116
rect 4668 3749 4811 4003
rect 4922 2154 5065 3749
rect 20799 3384 21037 3406
rect 6930 2154 13066 2197
rect 12760 1465 12998 1487
rect 3216 1340 3217 1366
<< metal1 >>
rect 1856 20837 11335 21274
rect 400 20400 2293 20837
rect 400 9565 836 20400
rect 1856 17575 2264 20197
rect 10898 20020 11335 20837
rect 16983 21212 17057 21786
rect 21755 21726 22025 21786
rect 22252 21726 22577 21786
rect 22749 21726 23129 21786
rect 23246 21726 23681 21786
rect 24159 21726 24521 21786
rect 24711 21726 25018 21786
rect 25263 21726 25514 21786
rect 25815 21726 26012 21786
rect 16983 20820 17108 21212
rect 20526 21018 20645 21092
rect 10303 19409 11191 19817
rect 20571 19437 20645 21018
rect 21755 20772 21815 21726
rect 22252 21026 22312 21726
rect 22749 21280 22809 21726
rect 23246 21534 23306 21726
rect 24461 21534 24521 21726
rect 22885 21474 23306 21534
rect 24460 21474 24881 21534
rect 24958 21280 25018 21726
rect 22388 21220 22809 21280
rect 24957 21220 25378 21280
rect 25455 21026 25515 21726
rect 21891 20966 22312 21026
rect 25454 20966 25875 21026
rect 25952 20772 26012 21726
rect 21394 20712 21815 20772
rect 25951 20712 26372 20772
rect 19345 19029 20645 19437
rect 20291 18017 20571 19029
rect 21926 18310 22362 20154
rect 21926 17873 22964 18310
rect 400 9128 1273 9565
rect 1476 9128 3474 9536
rect 836 1345 1273 9128
rect 836 908 2483 1345
rect 5009 1316 5417 2004
rect 13048 1624 13456 3923
rect 21087 3543 21495 9863
rect 22528 3340 22964 17873
rect 21058 2903 22964 3340
rect 21058 1421 21495 2903
rect 2686 1016 5417 1316
rect 13019 984 21495 1421
rect 13019 908 13456 984
rect 2046 472 13456 908
<< metal2 >>
rect 2294 20632 2502 20668
rect 2294 20496 2330 20632
rect 2466 20496 2502 20632
rect 2294 20460 2502 20496
rect 11336 20252 11544 20288
rect 11336 20116 11372 20252
rect 11508 20116 11544 20252
rect 11336 20080 11544 20116
rect 22138 17836 22346 17872
rect 1005 9738 1213 9774
rect 1005 9602 1041 9738
rect 1177 9602 1213 9738
rect 22138 17700 22174 17836
rect 22310 17700 22346 17836
rect 22138 17664 22346 17700
rect 1005 9566 1213 9602
rect 2215 1518 2423 1554
rect 2215 1382 2251 1518
rect 2387 1382 2423 1518
rect 20849 3244 21057 3280
rect 20849 3108 20885 3244
rect 21021 3108 21057 3244
rect 20849 3072 21057 3108
rect 2215 1346 2423 1382
rect 12810 1325 13018 1361
rect 12810 1189 12846 1325
rect 12982 1189 13018 1325
rect 12810 1153 13018 1189
<< via2 >>
rect 17126 21260 17182 21316
rect 17206 21260 17262 21316
rect 17286 21260 17342 21316
rect 17366 21260 17422 21316
rect 17446 21260 17502 21316
rect 17526 21260 17582 21316
rect 17606 21260 17662 21316
rect 17686 21260 17742 21316
rect 17766 21260 17822 21316
rect 17846 21260 17902 21316
rect 17926 21260 17982 21316
rect 18006 21260 18062 21316
rect 18086 21260 18142 21316
rect 18166 21260 18222 21316
rect 18246 21260 18302 21316
rect 18326 21260 18382 21316
rect 18406 21260 18462 21316
rect 18486 21260 18542 21316
rect 18566 21260 18622 21316
rect 18646 21260 18702 21316
rect 18726 21260 18782 21316
rect 18806 21260 18862 21316
rect 18886 21260 18942 21316
rect 18966 21260 19022 21316
rect 19046 21260 19102 21316
rect 19126 21260 19182 21316
rect 19206 21260 19262 21316
rect 19286 21260 19342 21316
rect 19366 21260 19422 21316
rect 19446 21260 19502 21316
rect 19526 21260 19582 21316
rect 19606 21260 19662 21316
rect 19686 21260 19742 21316
rect 19766 21260 19822 21316
rect 19846 21260 19902 21316
rect 19926 21260 19982 21316
rect 20006 21260 20062 21316
rect 20086 21260 20142 21316
rect 20166 21260 20222 21316
rect 20246 21260 20302 21316
rect 20326 21260 20382 21316
rect 20406 21260 20462 21316
rect 17126 20716 17182 20772
rect 17206 20716 17262 20772
rect 17286 20716 17342 20772
rect 17366 20716 17422 20772
rect 17446 20716 17502 20772
rect 17526 20716 17582 20772
rect 17606 20716 17662 20772
rect 17686 20716 17742 20772
rect 17766 20716 17822 20772
rect 17846 20716 17902 20772
rect 17926 20716 17982 20772
rect 18006 20716 18062 20772
rect 18086 20716 18142 20772
rect 18166 20716 18222 20772
rect 18246 20716 18302 20772
rect 18326 20716 18382 20772
rect 18406 20716 18462 20772
rect 18486 20716 18542 20772
rect 18566 20716 18622 20772
rect 18646 20716 18702 20772
rect 18726 20716 18782 20772
rect 18806 20716 18862 20772
rect 18886 20716 18942 20772
rect 18966 20716 19022 20772
rect 19046 20716 19102 20772
rect 19126 20716 19182 20772
rect 19206 20716 19262 20772
rect 19286 20716 19342 20772
rect 19366 20716 19422 20772
rect 19446 20716 19502 20772
rect 19526 20716 19582 20772
rect 19606 20716 19662 20772
rect 19686 20716 19742 20772
rect 19766 20716 19822 20772
rect 19846 20716 19902 20772
rect 19926 20716 19982 20772
rect 20006 20716 20062 20772
rect 20086 20716 20142 20772
rect 20166 20716 20222 20772
rect 20246 20716 20302 20772
rect 20326 20716 20382 20772
rect 20406 20716 20462 20772
rect 2330 20496 2466 20632
rect 21446 20405 21502 20461
rect 21536 20405 21592 20461
rect 21626 20405 21682 20461
rect 21716 20405 21772 20461
rect 21806 20405 21862 20461
rect 25953 20405 26009 20461
rect 26043 20405 26099 20461
rect 26133 20405 26189 20461
rect 26223 20405 26279 20461
rect 26313 20405 26369 20461
rect 11372 20116 11508 20252
rect 2366 18198 10262 18334
rect 11408 17818 19304 17954
rect 1041 9602 1177 9738
rect 3340 9638 3476 17534
rect 19875 9904 20011 17800
rect 22174 17700 22310 17836
rect 2251 1382 2387 1518
rect 4550 1418 4686 9314
rect 13089 5406 20985 5542
rect 5050 3488 12946 3624
rect 20885 3108 21021 3244
rect 12846 1189 12982 1325
<< metal3 >>
rect 0 22264 1938 22304
rect 0 10200 48 22264
rect 352 19724 1938 22264
rect 27746 22264 31464 22304
rect 2138 21808 16506 22085
rect 27746 21808 31112 22264
rect 2138 21316 31112 21808
rect 2138 21260 17126 21316
rect 17182 21260 17206 21316
rect 17262 21260 17286 21316
rect 17342 21260 17366 21316
rect 17422 21260 17446 21316
rect 17502 21260 17526 21316
rect 17582 21260 17606 21316
rect 17662 21260 17686 21316
rect 17742 21260 17766 21316
rect 17822 21260 17846 21316
rect 17902 21260 17926 21316
rect 17982 21260 18006 21316
rect 18062 21260 18086 21316
rect 18142 21260 18166 21316
rect 18222 21260 18246 21316
rect 18302 21260 18326 21316
rect 18382 21260 18406 21316
rect 18462 21260 18486 21316
rect 18542 21260 18566 21316
rect 18622 21260 18646 21316
rect 18702 21260 18726 21316
rect 18782 21260 18806 21316
rect 18862 21260 18886 21316
rect 18942 21260 18966 21316
rect 19022 21260 19046 21316
rect 19102 21260 19126 21316
rect 19182 21260 19206 21316
rect 19262 21260 19286 21316
rect 19342 21260 19366 21316
rect 19422 21260 19446 21316
rect 19502 21260 19526 21316
rect 19582 21260 19606 21316
rect 19662 21260 19686 21316
rect 19742 21260 19766 21316
rect 19822 21260 19846 21316
rect 19902 21260 19926 21316
rect 19982 21260 20006 21316
rect 20062 21260 20086 21316
rect 20142 21260 20166 21316
rect 20222 21260 20246 21316
rect 20302 21260 20326 21316
rect 20382 21260 20406 21316
rect 20462 21260 31112 21316
rect 2138 21116 31112 21260
rect 2138 20632 16734 21116
rect 2138 20496 2330 20632
rect 2466 20496 16734 20632
rect 2138 20252 16734 20496
rect 2138 20116 11372 20252
rect 11508 20116 16734 20252
rect 2138 19924 16734 20116
rect 16934 20772 22071 20916
rect 16934 20716 17126 20772
rect 17182 20716 17206 20772
rect 17262 20716 17286 20772
rect 17342 20716 17366 20772
rect 17422 20716 17446 20772
rect 17502 20716 17526 20772
rect 17582 20716 17606 20772
rect 17662 20716 17686 20772
rect 17742 20716 17766 20772
rect 17822 20716 17846 20772
rect 17902 20716 17926 20772
rect 17982 20716 18006 20772
rect 18062 20716 18086 20772
rect 18142 20716 18166 20772
rect 18222 20716 18246 20772
rect 18302 20716 18326 20772
rect 18382 20716 18406 20772
rect 18462 20716 18486 20772
rect 18542 20716 18566 20772
rect 18622 20716 18646 20772
rect 18702 20716 18726 20772
rect 18782 20716 18806 20772
rect 18862 20716 18886 20772
rect 18942 20716 18966 20772
rect 19022 20716 19046 20772
rect 19102 20716 19126 20772
rect 19182 20716 19206 20772
rect 19262 20716 19286 20772
rect 19342 20716 19366 20772
rect 19422 20716 19446 20772
rect 19502 20716 19526 20772
rect 19582 20716 19606 20772
rect 19662 20716 19686 20772
rect 19742 20716 19766 20772
rect 19822 20716 19846 20772
rect 19902 20716 19926 20772
rect 19982 20716 20006 20772
rect 20062 20716 20086 20772
rect 20142 20716 20166 20772
rect 20222 20716 20246 20772
rect 20302 20716 20326 20772
rect 20382 20716 20406 20772
rect 20462 20716 22071 20772
rect 16934 20461 22071 20716
rect 16934 20405 21446 20461
rect 21502 20405 21536 20461
rect 21592 20405 21626 20461
rect 21682 20405 21716 20461
rect 21772 20405 21806 20461
rect 21862 20405 22071 20461
rect 16934 19724 22071 20405
rect 352 18334 22071 19724
rect 352 18198 2366 18334
rect 10262 18228 22071 18334
rect 22271 20461 31112 21116
rect 22271 20405 25953 20461
rect 26009 20405 26043 20461
rect 26099 20405 26133 20461
rect 26189 20405 26223 20461
rect 26279 20405 26313 20461
rect 26369 20405 31112 20461
rect 10262 18198 21782 18228
rect 352 17954 21782 18198
rect 22271 18028 31112 20405
rect 352 17818 11408 17954
rect 19304 17818 21782 17954
rect 352 17800 21782 17818
rect 352 17534 19875 17800
rect 352 10200 3340 17534
rect 0 10130 3340 10200
rect 600 9738 2948 9930
rect 600 9602 1041 9738
rect 1177 9602 2948 9738
rect 600 9246 2948 9602
rect 3148 9638 3340 10130
rect 3476 9904 19875 17534
rect 20011 9904 21782 17800
rect 3476 9638 21782 9904
rect 3148 9446 21782 9638
rect 4358 9314 21782 9446
rect 600 1518 4158 9246
rect 600 1382 2251 1518
rect 2387 1382 4158 1518
rect 600 997 4158 1382
rect 4358 1418 4550 9314
rect 4686 5542 21782 9314
rect 4686 5406 13089 5542
rect 20985 5406 21782 5542
rect 4686 5214 21782 5406
rect 21982 17836 31112 18028
rect 21982 17700 22174 17836
rect 22310 17700 31112 17836
rect 4686 3624 20493 5214
rect 21982 5014 31112 17700
rect 4686 3488 5050 3624
rect 12946 3488 20493 3624
rect 4686 1717 20493 3488
rect 20693 3244 31112 5014
rect 20693 3108 20885 3244
rect 21021 3108 31112 3244
rect 4686 1418 12454 1717
rect 20693 1517 31112 3108
rect 4358 1226 12454 1418
rect 12654 1325 31112 1517
rect 12654 1189 12846 1325
rect 12982 1189 31112 1325
rect 12654 997 31112 1189
rect 600 40 31112 997
rect 31416 40 31464 22264
rect 600 0 31464 40
<< via3 >>
rect 48 10200 352 22264
rect 31112 40 31416 22264
<< metal4 >>
rect 0 22264 400 22304
rect 0 10200 48 22264
rect 352 10200 400 22264
rect 4294 22104 4354 22304
rect 4846 22104 4906 22304
rect 5398 22104 5458 22304
rect 5950 22104 6010 22304
rect 6502 22104 6562 22304
rect 7054 22104 7114 22304
rect 7606 22104 7666 22304
rect 8158 22104 8218 22304
rect 8710 22104 8770 22304
rect 9262 22104 9322 22304
rect 9814 22104 9874 22304
rect 10366 22104 10426 22304
rect 10918 22104 10978 22304
rect 11470 22104 11530 22304
rect 12022 22104 12082 22304
rect 12574 22104 12634 22304
rect 13126 22104 13186 22304
rect 13678 22104 13738 22304
rect 14230 22104 14290 22304
rect 14782 22104 14842 22304
rect 15334 22104 15394 22304
rect 15886 22104 15946 22304
rect 16438 22104 16498 22304
rect 16990 22104 17050 22304
rect 17542 22104 17602 22304
rect 18094 22104 18154 22304
rect 18646 22104 18706 22304
rect 19198 22104 19258 22304
rect 19750 22104 19810 22304
rect 20302 22104 20362 22304
rect 20854 22104 20914 22304
rect 21406 22104 21466 22304
rect 21958 22104 22018 22304
rect 22510 22104 22570 22304
rect 23062 22104 23122 22304
rect 23614 22104 23674 22304
rect 24166 22104 24226 22304
rect 24718 22104 24778 22304
rect 25270 22104 25330 22304
rect 25822 22104 25882 22304
rect 26374 22104 26434 22304
rect 26926 22104 26986 22304
rect 27478 22104 27538 22304
rect 31064 22264 31464 22304
rect 0 0 400 10200
rect 31064 40 31112 22264
rect 31416 40 31464 22264
rect 31064 0 31464 40
use dac_8bit  dac_8bit_0
timestamp 1699066547
transform 0 -1 26418 -1 0 21576
box 92 40 1432 5030
use driver  driver_0
timestamp 1699066547
transform -1 0 20538 0 -1 21336
box 0 0 3485 640
use inv_strvd  inv_strvd_0
timestamp 1699066547
transform 0 1 2220 1 0 1201
box 0 -1 8241 2591
use inv_strvd  inv_strvd_1
timestamp 1699066547
transform 1 0 2149 0 -1 20663
box 0 -1 8241 2591
use inv_strvd  inv_strvd_2
timestamp 1699066547
transform 1 0 11191 0 -1 20283
box 0 -1 8241 2591
use inv_strvd  inv_strvd_3
timestamp 1699066547
transform -1 0 13163 0 1 1158
box 0 -1 8241 2591
use inv_strvd  inv_strvd_4
timestamp 1699066547
transform 0 -1 22341 -1 0 18017
box 0 -1 8241 2591
use inv_strvd  inv_strvd_5
timestamp 1699066547
transform 0 1 1010 1 0 9421
box 0 -1 8241 2591
use inv_strvd  inv_strvd_6
timestamp 1699066547
transform -1 0 21202 0 1 3077
box 0 -1 8241 2591
use pin_connect  pin_connect_0
timestamp 1699066547
transform 1 0 27470 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_1
timestamp 1699066547
transform 1 0 26918 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_2
timestamp 1699066547
transform 1 0 26366 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_3
timestamp 1699066547
transform 1 0 25814 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_4
timestamp 1699066547
transform 1 0 25262 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_5
timestamp 1699066547
transform 1 0 24710 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_6
timestamp 1699066547
transform 1 0 24158 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_7
timestamp 1699066547
transform 1 0 23606 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_8
timestamp 1699066547
transform 1 0 23054 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_9
timestamp 1699066547
transform 1 0 22502 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_10
timestamp 1699066547
transform 1 0 21950 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_11
timestamp 1699066547
transform 1 0 21398 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_12
timestamp 1699066547
transform 1 0 20846 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_13
timestamp 1699066547
transform 1 0 20294 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_14
timestamp 1699066547
transform 1 0 19742 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_15
timestamp 1699066547
transform 1 0 19190 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_16
timestamp 1699066547
transform 1 0 18638 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_17
timestamp 1699066547
transform 1 0 18086 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_18
timestamp 1699066547
transform 1 0 17534 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_19
timestamp 1699066547
transform 1 0 16982 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_20
timestamp 1699066547
transform 1 0 16430 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_21
timestamp 1699066547
transform 1 0 15878 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_22
timestamp 1699066547
transform 1 0 15326 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_23
timestamp 1699066547
transform 1 0 14774 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_24
timestamp 1699066547
transform 1 0 14222 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_25
timestamp 1699066547
transform 1 0 13670 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_26
timestamp 1699066547
transform 1 0 13118 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_27
timestamp 1699066547
transform 1 0 12566 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_28
timestamp 1699066547
transform 1 0 12014 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_29
timestamp 1699066547
transform 1 0 11462 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_30
timestamp 1699066547
transform 1 0 10910 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_31
timestamp 1699066547
transform 1 0 10358 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_32
timestamp 1699066547
transform 1 0 9806 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_33
timestamp 1699066547
transform 1 0 9254 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_34
timestamp 1699066547
transform 1 0 8702 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_35
timestamp 1699066547
transform 1 0 8150 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_36
timestamp 1699066547
transform 1 0 7598 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_37
timestamp 1699066547
transform 1 0 7046 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_38
timestamp 1699066547
transform 1 0 6494 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_39
timestamp 1699066547
transform 1 0 5942 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_40
timestamp 1699066547
transform 1 0 5390 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_41
timestamp 1699066547
transform 1 0 4838 0 1 21786
box 0 0 76 518
use pin_connect  pin_connect_42
timestamp 1699066547
transform 1 0 4286 0 1 21786
box 0 0 76 518
use tt_um_template  tt_um_template_0
timestamp 1699066547
transform 1 0 0 0 1 0
box 0 0 1 1
<< labels >>
flabel metal4 s 31064 0 31464 22304 0 FreeSans 2000 0 0 0 VGND
port 2 nsew
rlabel metal4 s 26926 22104 26986 22304 4 clk
port 3 nsew
rlabel metal4 s 27478 22104 27538 22304 4 ena
port 4 nsew
rlabel metal4 s 26374 22104 26434 22304 4 rst_n
port 5 nsew
rlabel metal4 s 25822 22104 25882 22304 4 ui_in[0]
port 6 nsew
rlabel metal4 s 25270 22104 25330 22304 4 ui_in[1]
port 7 nsew
rlabel metal4 s 24718 22104 24778 22304 4 ui_in[2]
port 8 nsew
rlabel metal4 s 24166 22104 24226 22304 4 ui_in[3]
port 9 nsew
rlabel metal4 s 23614 22104 23674 22304 4 ui_in[4]
port 10 nsew
rlabel metal4 s 23062 22104 23122 22304 4 ui_in[5]
port 11 nsew
rlabel metal4 s 22510 22104 22570 22304 4 ui_in[6]
port 12 nsew
rlabel metal4 s 21958 22104 22018 22304 4 ui_in[7]
port 13 nsew
rlabel metal4 s 21406 22104 21466 22304 4 uio_in[0]
port 14 nsew
rlabel metal4 s 20854 22104 20914 22304 4 uio_in[1]
port 15 nsew
rlabel metal4 s 20302 22104 20362 22304 4 uio_in[2]
port 16 nsew
rlabel metal4 s 19750 22104 19810 22304 4 uio_in[3]
port 17 nsew
rlabel metal4 s 19198 22104 19258 22304 4 uio_in[4]
port 18 nsew
rlabel metal4 s 18646 22104 18706 22304 4 uio_in[5]
port 19 nsew
rlabel metal4 s 18094 22104 18154 22304 4 uio_in[6]
port 20 nsew
rlabel metal4 s 17542 22104 17602 22304 4 uio_in[7]
port 21 nsew
rlabel metal4 s 8158 22104 8218 22304 4 uio_oe[0]
port 22 nsew
rlabel metal4 s 7606 22104 7666 22304 4 uio_oe[1]
port 23 nsew
rlabel metal4 s 7054 22104 7114 22304 4 uio_oe[2]
port 24 nsew
rlabel metal4 s 6502 22104 6562 22304 4 uio_oe[3]
port 25 nsew
rlabel metal4 s 5950 22104 6010 22304 4 uio_oe[4]
port 26 nsew
rlabel metal4 s 5398 22104 5458 22304 4 uio_oe[5]
port 27 nsew
rlabel metal4 s 4846 22104 4906 22304 4 uio_oe[6]
port 28 nsew
rlabel metal4 s 4294 22104 4354 22304 4 uio_oe[7]
port 29 nsew
rlabel metal4 s 12574 22104 12634 22304 4 uio_out[0]
port 30 nsew
rlabel metal4 s 12022 22104 12082 22304 4 uio_out[1]
port 31 nsew
rlabel metal4 s 11470 22104 11530 22304 4 uio_out[2]
port 32 nsew
rlabel metal4 s 10918 22104 10978 22304 4 uio_out[3]
port 33 nsew
rlabel metal4 s 10366 22104 10426 22304 4 uio_out[4]
port 34 nsew
rlabel metal4 s 9814 22104 9874 22304 4 uio_out[5]
port 35 nsew
rlabel metal4 s 9262 22104 9322 22304 4 uio_out[6]
port 36 nsew
rlabel metal4 s 8710 22104 8770 22304 4 uio_out[7]
port 37 nsew
rlabel metal4 s 16990 22104 17050 22304 4 uo_out[0]
port 38 nsew
rlabel metal4 s 16438 22104 16498 22304 4 uo_out[1]
port 39 nsew
rlabel metal4 s 15886 22104 15946 22304 4 uo_out[2]
port 40 nsew
rlabel metal4 s 15334 22104 15394 22304 4 uo_out[3]
port 41 nsew
rlabel metal4 s 14782 22104 14842 22304 4 uo_out[4]
port 42 nsew
rlabel metal4 s 14230 22104 14290 22304 4 uo_out[5]
port 43 nsew
rlabel metal4 s 13678 22104 13738 22304 4 uo_out[6]
port 44 nsew
rlabel metal4 s 13126 22104 13186 22304 4 uo_out[7]
port 45 nsew
flabel metal4 s 0 0 400 22304 0 FreeSans 2000 0 0 0 VPWR
port 46 nsew
<< end >>
